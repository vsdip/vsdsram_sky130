magic
tech sky130A
timestamp 1617949095
<< nwell >>
rect 70 382 330 554
<< nmos >>
rect 123 159 138 285
rect 265 159 280 285
rect 146 110 188 125
rect 215 110 257 125
<< pmos >>
rect 123 400 138 455
rect 256 405 271 460
<< ndiff >>
rect 88 277 123 285
rect 88 260 96 277
rect 113 260 123 277
rect 88 184 123 260
rect 88 167 96 184
rect 113 167 123 184
rect 88 159 123 167
rect 138 277 188 285
rect 138 260 163 277
rect 180 260 188 277
rect 138 184 188 260
rect 138 167 163 184
rect 180 167 188 184
rect 138 159 188 167
rect 146 125 188 159
rect 215 277 265 285
rect 215 260 223 277
rect 240 260 265 277
rect 215 184 265 260
rect 215 167 223 184
rect 240 167 265 184
rect 215 159 265 167
rect 280 277 315 285
rect 280 260 290 277
rect 307 260 315 277
rect 280 184 315 260
rect 280 167 290 184
rect 307 167 315 184
rect 280 159 315 167
rect 215 125 257 159
rect 146 100 188 110
rect 146 83 163 100
rect 180 83 188 100
rect 146 76 188 83
rect 215 101 257 110
rect 215 84 223 101
rect 240 84 257 101
rect 215 76 257 84
<< pdiff >>
rect 88 447 123 455
rect 88 430 96 447
rect 113 430 123 447
rect 88 400 123 430
rect 138 425 173 455
rect 138 408 148 425
rect 165 408 173 425
rect 138 400 173 408
rect 221 452 256 460
rect 221 435 229 452
rect 246 435 256 452
rect 221 405 256 435
rect 271 430 306 460
rect 271 413 281 430
rect 298 413 306 430
rect 271 405 306 413
<< ndiffc >>
rect 96 260 113 277
rect 96 167 113 184
rect 163 260 180 277
rect 163 167 180 184
rect 223 260 240 277
rect 223 167 240 184
rect 290 260 307 277
rect 290 167 307 184
rect 163 83 180 100
rect 223 84 240 101
<< pdiffc >>
rect 96 430 113 447
rect 148 408 165 425
rect 229 435 246 452
rect 281 413 298 430
<< psubdiff >>
rect 80 61 118 73
rect 80 44 91 61
rect 108 44 118 61
rect 80 32 118 44
<< nsubdiff >>
rect 88 508 141 535
rect 88 491 100 508
rect 117 491 141 508
rect 88 482 141 491
<< psubdiffcont >>
rect 91 44 108 61
<< nsubdiffcont >>
rect 100 491 117 508
<< poly >>
rect 123 455 138 468
rect 256 460 271 473
rect 123 389 138 400
rect 123 381 235 389
rect 123 374 210 381
rect 123 285 138 374
rect 202 364 210 374
rect 227 364 235 381
rect 202 356 235 364
rect 160 327 193 335
rect 160 310 168 327
rect 185 324 193 327
rect 256 324 271 405
rect 185 310 280 324
rect 160 309 280 310
rect 160 302 193 309
rect 265 285 280 309
rect 123 146 138 159
rect 265 146 280 159
rect 70 117 146 125
rect 70 110 96 117
rect 88 100 96 110
rect 113 110 146 117
rect 188 110 215 125
rect 257 110 330 125
rect 113 100 121 110
rect 88 92 121 100
<< polycont >>
rect 210 364 227 381
rect 168 310 185 327
rect 96 100 113 117
<< locali >>
rect 92 508 125 516
rect 92 491 100 508
rect 117 491 125 508
rect 92 483 125 491
rect 213 509 245 517
rect 213 492 220 509
rect 237 492 245 509
rect 213 484 245 492
rect 274 508 306 516
rect 274 491 281 508
rect 298 491 306 508
rect 98 455 115 483
rect 221 460 238 484
rect 274 483 306 491
rect 88 447 121 455
rect 88 430 96 447
rect 113 430 121 447
rect 221 452 254 460
rect 221 435 229 452
rect 246 435 254 452
rect 281 438 298 483
rect 88 422 121 430
rect 140 425 173 433
rect 140 408 148 425
rect 165 408 173 425
rect 140 400 173 408
rect 221 427 254 435
rect 273 430 306 438
rect 155 335 172 400
rect 221 389 238 427
rect 273 413 281 430
rect 298 413 306 430
rect 273 405 306 413
rect 202 381 238 389
rect 202 364 210 381
rect 227 364 238 381
rect 202 356 238 364
rect 155 327 193 335
rect 155 310 168 327
rect 185 310 193 327
rect 155 302 193 310
rect 155 285 172 302
rect 221 285 238 356
rect 88 277 121 285
rect 88 260 96 277
rect 113 260 121 277
rect 88 231 121 260
rect 155 277 188 285
rect 155 260 163 277
rect 180 260 188 277
rect 155 252 188 260
rect 215 277 248 285
rect 215 260 223 277
rect 240 260 248 277
rect 215 252 248 260
rect 282 277 315 285
rect 282 260 290 277
rect 307 260 315 277
rect 282 231 315 260
rect 88 214 315 231
rect 88 184 121 214
rect 88 167 96 184
rect 113 167 121 184
rect 88 159 121 167
rect 155 184 188 192
rect 155 167 163 184
rect 180 167 188 184
rect 155 159 188 167
rect 215 184 248 192
rect 215 167 223 184
rect 240 167 248 184
rect 215 159 248 167
rect 282 184 315 214
rect 282 167 290 184
rect 307 167 315 184
rect 282 159 315 167
rect 88 117 121 125
rect 88 100 96 117
rect 113 100 121 117
rect 88 92 121 100
rect 155 100 188 108
rect 155 83 163 100
rect 180 83 188 100
rect 155 76 188 83
rect 215 101 248 109
rect 215 84 223 101
rect 240 84 248 101
rect 215 76 248 84
rect 164 69 181 76
rect 83 61 116 69
rect 83 44 91 61
rect 108 44 116 61
rect 215 69 232 76
rect 298 55 315 159
rect 83 35 116 44
rect 298 30 315 38
<< viali >>
rect 100 491 117 508
rect 220 492 237 509
rect 281 491 298 508
rect 210 364 227 381
rect 168 310 185 327
rect 96 100 113 117
rect 91 44 108 61
rect 164 52 181 69
rect 215 52 232 69
rect 298 38 315 55
<< metal1 >>
rect 0 509 400 554
rect 92 508 125 509
rect 92 491 100 508
rect 117 491 125 508
rect 92 483 125 491
rect 213 492 220 509
rect 237 492 245 509
rect 213 484 245 492
rect 274 508 306 509
rect 274 491 281 508
rect 298 491 306 508
rect 274 483 306 491
rect 204 381 233 387
rect 204 364 210 381
rect 227 364 233 381
rect 204 358 233 364
rect 162 327 191 333
rect 162 310 168 327
rect 185 310 191 327
rect 162 304 191 310
rect 90 117 119 123
rect 90 107 96 117
rect 88 100 96 107
rect 113 107 119 117
rect 113 100 121 107
rect 88 92 121 100
rect 156 73 188 76
rect 85 61 114 68
rect 85 44 91 61
rect 108 44 114 61
rect 156 47 159 73
rect 185 47 188 73
rect 156 44 188 47
rect 207 73 239 76
rect 207 47 210 73
rect 236 47 239 73
rect 207 44 239 47
rect 290 55 320 62
rect 85 21 114 44
rect 290 38 298 55
rect 315 38 320 55
rect 290 21 320 38
rect 0 -20 400 21
<< via1 >>
rect 159 69 185 73
rect 159 52 164 69
rect 164 52 181 69
rect 181 52 185 69
rect 159 47 185 52
rect 210 69 236 73
rect 210 52 215 69
rect 215 52 232 69
rect 232 52 236 69
rect 210 47 236 52
<< metal2 >>
rect 123 65 137 554
rect 156 73 188 76
rect 156 65 159 73
rect 123 51 159 65
rect 123 -20 137 51
rect 156 47 159 51
rect 185 47 188 73
rect 156 44 188 47
rect 207 73 239 76
rect 207 47 210 73
rect 236 66 239 73
rect 265 66 279 554
rect 236 52 279 66
rect 236 47 239 52
rect 207 44 239 47
rect 265 -20 279 52
<< labels >>
flabel locali s 213 367 224 378 0 FreeSans 200 0 0 0 qb
port 10 nsew
flabel metal2 s 265 52 278 66 0 FreeSans 200 0 0 0 br
port 16 nsew
flabel metal2 s 123 51 136 65 0 FreeSans 200 0 0 0 bl
port 17 nsew
flabel metal1 s 98 102 109 113 0 FreeSans 200 0 0 0 wl
port 5 nsew
flabel metal1 s 257 -5 268 6 0 FreeSans 200 0 0 0 gnd
port 3 nsew
flabel metal1 s 181 520 223 540 0 FreeSans 200 0 0 0 vdd
port 1 nsew
flabel locali s 172 314 183 325 0 FreeSans 200 0 0 0 q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 400 532
<< end >>
