magic
tech sky130A
timestamp 1617954257
<< nwell >>
rect 0 281 1313 461
<< nmos >>
rect 81 85 96 127
rect 224 85 239 127
rect 345 85 360 127
rect 516 85 531 127
rect 611 85 626 127
rect 804 85 819 127
rect 925 85 940 127
rect 1120 85 1135 127
rect 1215 85 1230 127
<< pmos >>
rect 81 299 96 354
rect 224 299 239 354
rect 345 299 360 354
rect 516 299 531 354
rect 611 299 626 354
rect 804 299 819 354
rect 925 299 940 354
rect 1120 299 1135 354
rect 1215 299 1230 354
<< ndiff >>
rect 35 116 81 127
rect 35 99 45 116
rect 62 99 81 116
rect 35 85 81 99
rect 96 116 142 127
rect 96 99 114 116
rect 131 99 142 116
rect 96 85 142 99
rect 178 116 224 127
rect 178 99 188 116
rect 205 99 224 116
rect 178 85 224 99
rect 239 116 345 127
rect 239 99 298 116
rect 315 99 345 116
rect 239 85 345 99
rect 360 116 428 127
rect 360 99 393 116
rect 410 99 428 116
rect 360 85 428 99
rect 463 115 516 127
rect 463 98 476 115
rect 493 98 516 115
rect 463 85 516 98
rect 531 116 611 127
rect 531 99 564 116
rect 581 99 611 116
rect 531 85 611 99
rect 626 116 688 127
rect 626 99 639 116
rect 656 99 688 116
rect 626 85 688 99
rect 739 116 804 127
rect 739 99 768 116
rect 785 99 804 116
rect 739 85 804 99
rect 819 116 925 127
rect 819 99 878 116
rect 895 99 925 116
rect 819 85 925 99
rect 940 116 1019 127
rect 940 99 973 116
rect 990 99 1019 116
rect 940 85 1019 99
rect 1064 116 1120 127
rect 1064 99 1080 116
rect 1097 99 1120 116
rect 1064 85 1120 99
rect 1135 116 1215 127
rect 1135 99 1168 116
rect 1185 99 1215 116
rect 1135 85 1215 99
rect 1230 116 1270 127
rect 1230 99 1243 116
rect 1260 99 1270 116
rect 1230 85 1270 99
<< pdiff >>
rect 35 336 81 354
rect 35 319 45 336
rect 62 319 81 336
rect 35 299 81 319
rect 96 336 142 354
rect 96 319 114 336
rect 131 319 142 336
rect 96 299 142 319
rect 178 336 224 354
rect 178 319 188 336
rect 205 319 224 336
rect 178 299 224 319
rect 239 336 345 354
rect 239 319 298 336
rect 315 319 345 336
rect 239 299 345 319
rect 360 336 428 354
rect 360 319 393 336
rect 410 319 428 336
rect 360 299 428 319
rect 463 336 516 354
rect 463 319 481 336
rect 498 319 516 336
rect 463 299 516 319
rect 531 336 611 354
rect 531 319 564 336
rect 581 319 611 336
rect 531 299 611 319
rect 626 336 689 354
rect 626 319 639 336
rect 656 319 689 336
rect 626 299 689 319
rect 740 336 804 354
rect 740 319 768 336
rect 785 319 804 336
rect 740 299 804 319
rect 819 336 925 354
rect 819 319 878 336
rect 895 319 925 336
rect 819 299 925 319
rect 940 336 1019 354
rect 940 319 973 336
rect 990 319 1019 336
rect 940 299 1019 319
rect 1064 336 1120 354
rect 1064 319 1077 336
rect 1094 319 1120 336
rect 1064 299 1120 319
rect 1135 336 1215 354
rect 1135 319 1168 336
rect 1185 319 1215 336
rect 1135 299 1215 319
rect 1230 336 1270 354
rect 1230 319 1243 336
rect 1260 319 1270 336
rect 1230 299 1270 319
<< ndiffc >>
rect 45 99 62 116
rect 114 99 131 116
rect 188 99 205 116
rect 298 99 315 116
rect 393 99 410 116
rect 476 98 493 115
rect 564 99 581 116
rect 639 99 656 116
rect 768 99 785 116
rect 878 99 895 116
rect 973 99 990 116
rect 1080 99 1097 116
rect 1168 99 1185 116
rect 1243 99 1260 116
<< pdiffc >>
rect 45 319 62 336
rect 114 319 131 336
rect 188 319 205 336
rect 298 319 315 336
rect 393 319 410 336
rect 481 319 498 336
rect 564 319 581 336
rect 639 319 656 336
rect 768 319 785 336
rect 878 319 895 336
rect 973 319 990 336
rect 1077 319 1094 336
rect 1168 319 1185 336
rect 1243 319 1260 336
<< psubdiff >>
rect 163 51 204 58
rect 163 34 175 51
rect 192 34 204 51
rect 163 -14 204 34
rect 267 51 308 58
rect 267 34 279 51
rect 296 34 308 51
rect 267 -14 308 34
rect 378 51 419 58
rect 378 34 390 51
rect 407 34 419 51
rect 378 -14 419 34
rect 743 51 784 58
rect 743 34 755 51
rect 772 34 784 51
rect 743 -14 784 34
rect 847 51 888 58
rect 847 34 859 51
rect 876 34 888 51
rect 847 -14 888 34
rect 958 51 999 58
rect 958 34 970 51
rect 987 34 999 51
rect 958 -14 999 34
rect 1068 51 1109 58
rect 1068 34 1080 51
rect 1097 34 1109 51
rect 1068 -14 1109 34
<< nsubdiff >>
rect 178 407 231 443
rect 178 390 195 407
rect 212 390 231 407
rect 178 381 231 390
rect 330 407 383 443
rect 330 390 347 407
rect 364 390 383 407
rect 330 381 383 390
rect 482 407 535 443
rect 482 390 499 407
rect 516 390 535 407
rect 482 381 535 390
rect 758 407 811 443
rect 758 390 775 407
rect 792 390 811 407
rect 758 381 811 390
rect 910 407 963 443
rect 910 390 927 407
rect 944 390 963 407
rect 910 381 963 390
rect 1087 407 1140 443
rect 1087 390 1104 407
rect 1121 390 1140 407
rect 1087 381 1140 390
rect 1222 407 1275 443
rect 1222 390 1239 407
rect 1256 390 1275 407
rect 1222 381 1275 390
<< psubdiffcont >>
rect 175 34 192 51
rect 279 34 296 51
rect 390 34 407 51
rect 755 34 772 51
rect 859 34 876 51
rect 970 34 987 51
rect 1080 34 1097 51
<< nsubdiffcont >>
rect 195 390 212 407
rect 347 390 364 407
rect 499 390 516 407
rect 775 390 792 407
rect 927 390 944 407
rect 1104 390 1121 407
rect 1239 390 1256 407
<< poly >>
rect 81 354 96 369
rect 224 354 239 369
rect 345 354 360 369
rect 516 354 531 369
rect 611 354 626 369
rect 804 354 819 369
rect 925 354 940 369
rect 1120 354 1135 369
rect 1215 354 1230 369
rect 81 227 96 299
rect 224 227 239 299
rect 345 277 360 299
rect 516 279 531 299
rect 336 269 369 277
rect 336 252 344 269
rect 361 252 369 269
rect 336 244 369 252
rect 516 271 549 279
rect 516 254 524 271
rect 541 254 549 271
rect 516 246 549 254
rect 81 223 239 227
rect 81 215 369 223
rect 81 207 344 215
rect 25 183 58 187
rect 81 183 96 207
rect 336 198 344 207
rect 361 198 369 215
rect 336 190 369 198
rect 25 179 96 183
rect 25 162 33 179
rect 50 168 96 179
rect 50 162 58 168
rect 25 154 58 162
rect 81 127 96 168
rect 224 175 257 183
rect 224 158 232 175
rect 249 158 257 175
rect 224 150 257 158
rect 224 127 239 150
rect 345 127 360 190
rect 516 127 531 246
rect 611 177 626 299
rect 744 270 777 277
rect 804 270 819 299
rect 925 277 940 299
rect 744 269 819 270
rect 744 252 752 269
rect 769 255 819 269
rect 769 252 777 255
rect 744 244 777 252
rect 804 223 819 255
rect 916 269 949 277
rect 916 252 924 269
rect 941 252 949 269
rect 916 244 949 252
rect 1120 242 1135 299
rect 1120 234 1153 242
rect 804 215 949 223
rect 804 207 924 215
rect 916 198 924 207
rect 941 198 949 215
rect 916 190 949 198
rect 1120 217 1128 234
rect 1145 217 1153 234
rect 1120 209 1153 217
rect 593 169 626 177
rect 593 152 601 169
rect 618 152 626 169
rect 593 144 626 152
rect 611 127 626 144
rect 804 171 837 179
rect 804 154 812 171
rect 829 154 837 171
rect 804 146 837 154
rect 804 127 819 146
rect 925 127 940 190
rect 1120 127 1135 209
rect 1215 178 1230 299
rect 1197 170 1230 178
rect 1197 153 1205 170
rect 1222 153 1230 170
rect 1197 145 1230 153
rect 1215 127 1230 145
rect 81 70 96 85
rect 224 70 239 85
rect 345 70 360 85
rect 516 70 531 85
rect 611 70 626 85
rect 804 70 819 85
rect 925 70 940 85
rect 1120 70 1135 85
rect 1215 70 1230 85
<< polycont >>
rect 344 252 361 269
rect 524 254 541 271
rect 344 198 361 215
rect 33 162 50 179
rect 232 158 249 175
rect 752 252 769 269
rect 924 252 941 269
rect 924 198 941 215
rect 1128 217 1145 234
rect 601 152 618 169
rect 812 154 829 171
rect 1205 153 1222 170
<< locali >>
rect 0 410 1313 443
rect 43 344 63 410
rect 178 407 231 410
rect 178 390 195 407
rect 212 390 231 407
rect 178 381 231 390
rect 330 407 383 410
rect 330 390 347 407
rect 364 390 383 407
rect 330 381 383 390
rect 482 407 535 410
rect 482 390 499 407
rect 516 390 535 407
rect 482 381 535 390
rect 559 344 579 410
rect 758 407 811 410
rect 758 390 775 407
rect 792 390 811 407
rect 758 381 811 390
rect 910 407 963 410
rect 910 390 927 407
rect 944 390 963 407
rect 910 381 963 390
rect 1087 407 1140 410
rect 1087 390 1104 407
rect 1121 390 1140 407
rect 1087 381 1140 390
rect 1163 344 1183 410
rect 1222 407 1275 410
rect 1222 390 1239 407
rect 1256 390 1275 407
rect 1222 381 1275 390
rect 37 336 70 344
rect 37 319 45 336
rect 62 319 70 336
rect 37 311 70 319
rect 106 336 139 344
rect 106 319 114 336
rect 131 319 139 336
rect 106 311 139 319
rect 180 336 213 344
rect 180 319 188 336
rect 205 319 213 336
rect 180 311 213 319
rect 290 336 323 344
rect 290 319 298 336
rect 315 319 323 336
rect 290 311 323 319
rect 385 340 418 344
rect 473 340 506 344
rect 385 336 506 340
rect 385 319 393 336
rect 410 319 481 336
rect 498 319 506 336
rect 385 315 506 319
rect 385 311 418 315
rect 473 311 506 315
rect 556 336 589 344
rect 556 319 564 336
rect 581 319 589 336
rect 556 311 589 319
rect 631 336 793 344
rect 631 319 639 336
rect 656 319 768 336
rect 785 319 793 336
rect 631 311 793 319
rect 870 336 903 344
rect 870 319 878 336
rect 895 319 903 336
rect 870 311 903 319
rect 965 336 998 344
rect 965 319 973 336
rect 990 335 998 336
rect 1069 336 1102 344
rect 1069 335 1077 336
rect 990 319 1077 335
rect 1094 319 1102 336
rect 965 315 1102 319
rect 965 311 998 315
rect 1069 311 1102 315
rect 1160 336 1193 344
rect 1160 319 1168 336
rect 1185 319 1193 336
rect 1160 311 1193 319
rect 1235 336 1268 344
rect 1235 319 1243 336
rect 1260 319 1268 336
rect 1235 311 1268 319
rect 25 179 58 187
rect 113 181 133 311
rect 180 308 203 311
rect 175 302 203 308
rect 175 285 180 302
rect 197 285 203 302
rect 175 280 203 285
rect 25 161 33 179
rect 50 161 58 179
rect 25 154 58 161
rect 112 175 141 181
rect 112 158 118 175
rect 135 158 141 175
rect 112 152 141 158
rect 113 124 133 152
rect 183 124 203 280
rect 224 175 257 183
rect 295 181 315 311
rect 336 269 369 277
rect 336 252 344 269
rect 361 252 369 269
rect 336 244 369 252
rect 336 215 369 223
rect 336 198 344 215
rect 361 198 369 215
rect 336 190 369 198
rect 224 158 232 175
rect 249 158 257 175
rect 224 150 257 158
rect 283 173 315 181
rect 283 156 289 173
rect 306 156 315 173
rect 283 150 315 156
rect 295 124 315 150
rect 390 124 410 311
rect 516 272 549 279
rect 644 272 664 311
rect 516 271 664 272
rect 516 254 524 271
rect 541 254 664 271
rect 516 252 664 254
rect 516 246 549 252
rect 593 169 626 177
rect 593 152 601 169
rect 618 152 626 169
rect 593 144 626 152
rect 644 124 664 252
rect 744 269 777 277
rect 744 252 752 269
rect 769 252 777 269
rect 744 244 777 252
rect 875 179 895 311
rect 916 269 949 277
rect 916 252 924 269
rect 941 252 949 269
rect 916 244 949 252
rect 916 215 949 223
rect 916 198 924 215
rect 941 198 949 215
rect 916 190 949 198
rect 804 171 837 179
rect 804 154 812 171
rect 829 154 837 171
rect 804 146 837 154
rect 863 171 895 179
rect 863 154 869 171
rect 886 154 895 171
rect 863 148 895 154
rect 875 124 895 148
rect 970 124 990 311
rect 1062 235 1153 242
rect 1248 235 1268 311
rect 1062 234 1268 235
rect 1062 217 1069 234
rect 1086 217 1128 234
rect 1145 217 1268 234
rect 1062 215 1268 217
rect 1062 210 1153 215
rect 1120 209 1153 210
rect 1197 170 1230 178
rect 1197 153 1205 170
rect 1222 153 1230 170
rect 1197 145 1230 153
rect 1248 124 1268 215
rect 37 116 70 124
rect 37 99 45 116
rect 62 99 70 116
rect 37 91 70 99
rect 106 116 139 124
rect 106 99 114 116
rect 131 99 139 116
rect 106 91 139 99
rect 180 116 213 124
rect 180 99 188 116
rect 205 99 213 116
rect 180 91 213 99
rect 290 116 323 124
rect 290 99 298 116
rect 315 99 323 116
rect 290 91 323 99
rect 385 116 418 124
rect 385 99 393 116
rect 410 115 418 116
rect 468 115 501 123
rect 410 99 476 115
rect 385 98 476 99
rect 493 98 501 115
rect 385 95 501 98
rect 385 91 418 95
rect 43 17 63 91
rect 468 90 501 95
rect 556 116 589 124
rect 556 99 564 116
rect 581 99 589 116
rect 556 91 589 99
rect 163 51 204 58
rect 163 34 175 51
rect 192 34 204 51
rect 163 17 204 34
rect 267 51 308 58
rect 267 34 279 51
rect 296 34 308 51
rect 267 17 308 34
rect 378 51 419 58
rect 378 34 390 51
rect 407 34 419 51
rect 378 17 419 34
rect 569 17 589 91
rect 631 116 793 124
rect 631 99 639 116
rect 656 99 768 116
rect 785 99 793 116
rect 631 90 793 99
rect 870 116 903 124
rect 870 99 878 116
rect 895 99 903 116
rect 870 91 903 99
rect 965 116 998 124
rect 965 99 973 116
rect 990 115 998 116
rect 1072 116 1105 124
rect 1072 115 1080 116
rect 990 99 1080 115
rect 1097 99 1105 116
rect 965 95 1105 99
rect 965 91 998 95
rect 1072 91 1105 95
rect 1160 116 1193 124
rect 1160 99 1168 116
rect 1185 99 1193 116
rect 1160 91 1193 99
rect 1235 116 1268 124
rect 1235 99 1243 116
rect 1260 99 1268 116
rect 1235 91 1268 99
rect 743 51 784 58
rect 743 34 755 51
rect 772 34 784 51
rect 743 17 784 34
rect 847 51 888 58
rect 847 34 859 51
rect 876 34 888 51
rect 847 17 888 34
rect 958 51 999 58
rect 958 34 970 51
rect 987 34 999 51
rect 958 17 999 34
rect 1068 51 1109 58
rect 1068 34 1080 51
rect 1097 34 1109 51
rect 1068 17 1109 34
rect 1173 17 1193 91
rect 0 -14 1313 17
<< viali >>
rect 195 390 212 407
rect 347 390 364 407
rect 499 390 516 407
rect 775 390 792 407
rect 927 390 944 407
rect 1104 390 1121 407
rect 1239 390 1256 407
rect 180 285 197 302
rect 33 162 50 178
rect 33 161 50 162
rect 118 158 135 175
rect 344 252 361 269
rect 344 198 361 215
rect 232 158 249 175
rect 289 156 306 173
rect 601 152 618 169
rect 752 252 769 269
rect 924 252 941 269
rect 812 154 829 171
rect 869 154 886 171
rect 1069 217 1086 234
rect 1205 153 1222 170
rect 175 34 192 51
rect 279 34 296 51
rect 390 34 407 51
rect 755 34 772 51
rect 859 34 876 51
rect 970 34 987 51
rect 1080 34 1097 51
<< metal1 >>
rect 0 407 1313 449
rect 0 404 195 407
rect 178 390 195 404
rect 212 404 347 407
rect 212 390 231 404
rect 178 381 231 390
rect 330 390 347 404
rect 364 404 499 407
rect 364 390 383 404
rect 330 381 383 390
rect 482 390 499 404
rect 516 404 775 407
rect 516 390 535 404
rect 482 381 535 390
rect 758 390 775 404
rect 792 404 927 407
rect 792 390 811 404
rect 758 381 811 390
rect 910 390 927 404
rect 944 404 1104 407
rect 944 390 963 404
rect 910 381 963 390
rect 1087 390 1104 404
rect 1121 404 1239 407
rect 1121 390 1140 404
rect 1087 381 1140 390
rect 1222 390 1239 404
rect 1256 404 1313 407
rect 1256 390 1275 404
rect 1222 381 1275 390
rect 174 307 208 310
rect 174 281 178 307
rect 204 281 208 307
rect 174 278 208 281
rect 336 269 369 277
rect 336 265 344 269
rect 228 252 344 265
rect 361 265 369 269
rect 744 269 777 277
rect 744 265 752 269
rect 361 252 752 265
rect 769 252 777 269
rect 916 269 949 277
rect 916 265 924 269
rect 228 245 777 252
rect 25 183 56 186
rect 228 183 248 245
rect 336 244 369 245
rect 744 244 777 245
rect 808 252 924 265
rect 941 252 949 269
rect 808 245 949 252
rect 336 220 369 223
rect 808 220 828 245
rect 916 244 949 245
rect 336 215 828 220
rect 336 198 344 215
rect 361 198 828 215
rect 1030 239 1093 242
rect 1030 213 1033 239
rect 1059 234 1093 239
rect 1059 217 1069 234
rect 1086 217 1093 234
rect 1059 213 1093 217
rect 1030 210 1093 213
rect 336 195 828 198
rect 336 190 369 195
rect 25 157 27 183
rect 53 157 56 183
rect 25 154 56 157
rect 112 175 141 181
rect 224 175 257 183
rect 112 158 118 175
rect 135 158 232 175
rect 249 158 257 175
rect 112 155 257 158
rect 112 152 141 155
rect 224 150 257 155
rect 283 175 313 181
rect 808 179 828 195
rect 593 175 626 177
rect 283 173 626 175
rect 283 156 289 173
rect 306 169 626 173
rect 306 156 601 169
rect 283 154 601 156
rect 283 150 313 154
rect 593 152 601 154
rect 618 152 626 169
rect 593 144 626 152
rect 804 171 837 179
rect 804 154 812 171
rect 829 154 837 171
rect 804 146 837 154
rect 863 175 893 179
rect 1196 175 1230 178
rect 863 171 1230 175
rect 863 154 869 171
rect 886 170 1230 171
rect 886 155 1205 170
rect 886 154 893 155
rect 863 148 893 154
rect 1196 153 1205 155
rect 1222 153 1230 170
rect 1196 145 1230 153
rect 163 51 204 58
rect 163 34 175 51
rect 192 34 204 51
rect 163 21 204 34
rect 267 51 308 58
rect 267 34 279 51
rect 296 34 308 51
rect 267 21 308 34
rect 378 51 419 58
rect 378 34 390 51
rect 407 34 419 51
rect 378 21 419 34
rect 743 51 784 58
rect 743 34 755 51
rect 772 34 784 51
rect 743 21 784 34
rect 847 51 888 58
rect 847 34 859 51
rect 876 34 888 51
rect 847 21 888 34
rect 958 51 999 58
rect 958 34 970 51
rect 987 34 999 51
rect 958 21 999 34
rect 1068 51 1109 58
rect 1068 34 1080 51
rect 1097 34 1109 51
rect 1068 21 1109 34
rect 0 -20 1313 21
<< via1 >>
rect 178 302 204 307
rect 178 285 180 302
rect 180 285 197 302
rect 197 285 204 302
rect 178 281 204 285
rect 1033 213 1059 239
rect 27 178 53 183
rect 27 161 33 178
rect 33 161 50 178
rect 50 161 53 178
rect 27 157 53 161
<< metal2 >>
rect 174 307 208 310
rect 174 281 178 307
rect 204 281 208 307
rect 174 278 208 281
rect 1030 239 1062 242
rect 1030 213 1033 239
rect 1059 213 1062 239
rect 1030 210 1062 213
rect 25 183 56 186
rect 25 157 27 183
rect 53 157 56 183
rect 25 154 56 157
<< labels >>
flabel locali s 975 320 985 332 0 FreeSans 200 0 0 0 net5
flabel metal2 s 1033 213 1059 239 0 FreeSans 400 0 0 0 Q
port 9 nsew
flabel metal2 s 178 281 204 307 0 FreeSans 400 0 0 0 D
port 2 nsew
flabel metal1 s 609 416 648 436 0 FreeSans 400 0 0 0 vdd
port 0 nsew
flabel locali s 396 190 404 198 0 FreeSans 200 0 0 0 net2
flabel locali s 652 158 660 166 0 FreeSans 200 0 0 0 net3
flabel locali s 234 159 245 172 0 FreeSans 240 0 0 0 clkb
flabel metal1 s 556 1 691 34 0 FreeSans 400 0 0 0 gnd
port 1 nsew
flabel locali s 292 160 300 167 0 FreeSans 200 0 0 0 net1
flabel locali s 874 157 882 164 0 FreeSans 200 0 0 0 net4
flabel metal2 s 27 157 53 183 0 FreeSans 240 0 0 0 clk
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1313 426
<< end >>
