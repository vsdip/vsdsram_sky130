VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130A
   CLASS BLOCK ;
   SIZE 72.96 BY 127.7 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  13.91 -11.08 14.65 -10.34 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  27.0 -11.08 27.74 -10.34 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -14.65 126.96 -13.91 127.7 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -11.08 126.96 -10.34 127.7 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.46 126.96 -12.72 127.7 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -12.27 126.96 -11.53 127.7 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -53.92 -7.51 -53.18 -6.77 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -50.35 -11.08 -49.61 -10.34 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -21.79 -11.08 -21.05 -10.34 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  72.22 16.29 72.96 17.03 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  72.22 11.53 72.96 12.27 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -53.92 -6.32 -51.99 -4.39 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -53.92 -11.08 -51.99 -9.15 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  54.89 40.95 58.89 41.4 ;
      RECT  54.89 35.66 58.89 36.07 ;
      RECT  55.77 36.78 56.1 36.93 ;
      RECT  57.79 36.07 58.09 36.48 ;
      RECT  55.79 36.93 56.08 37.09 ;
      RECT  55.74 36.07 56.03 36.54 ;
      RECT  56.45 36.3 56.77 36.62 ;
      RECT  57.63 40.69 57.95 40.95 ;
      RECT  56.51 38.9 56.8 39.19 ;
      RECT  56.96 36.3 57.28 36.62 ;
      RECT  56.93 39.44 57.22 39.73 ;
      RECT  55.81 40.69 56.14 40.95 ;
      RECT  54.89 41.41 58.89 40.96 ;
      RECT  54.89 46.7 58.89 46.29 ;
      RECT  55.77 45.58 56.1 45.43 ;
      RECT  57.79 46.29 58.09 45.88 ;
      RECT  55.79 45.43 56.08 45.27 ;
      RECT  55.74 46.29 56.03 45.82 ;
      RECT  56.45 46.06 56.77 45.74 ;
      RECT  57.63 41.67 57.95 41.41 ;
      RECT  56.51 43.46 56.8 43.17 ;
      RECT  56.96 46.06 57.28 45.74 ;
      RECT  56.93 42.92 57.22 42.63 ;
      RECT  55.81 41.67 56.14 41.41 ;
      RECT  54.89 51.59 58.89 52.04 ;
      RECT  54.89 46.3 58.89 46.71 ;
      RECT  55.77 47.42 56.1 47.57 ;
      RECT  57.79 46.71 58.09 47.12 ;
      RECT  55.79 47.57 56.08 47.73 ;
      RECT  55.74 46.71 56.03 47.18 ;
      RECT  56.45 46.94 56.77 47.26 ;
      RECT  57.63 51.33 57.95 51.59 ;
      RECT  56.51 49.54 56.8 49.83 ;
      RECT  56.96 46.94 57.28 47.26 ;
      RECT  56.93 50.08 57.22 50.37 ;
      RECT  55.81 51.33 56.14 51.59 ;
      RECT  54.89 52.05 58.89 51.6 ;
      RECT  54.89 57.34 58.89 56.93 ;
      RECT  55.77 56.22 56.1 56.07 ;
      RECT  57.79 56.93 58.09 56.52 ;
      RECT  55.79 56.07 56.08 55.91 ;
      RECT  55.74 56.93 56.03 56.46 ;
      RECT  56.45 56.7 56.77 56.38 ;
      RECT  57.63 52.31 57.95 52.05 ;
      RECT  56.51 54.1 56.8 53.81 ;
      RECT  56.96 56.7 57.28 56.38 ;
      RECT  56.93 53.56 57.22 53.27 ;
      RECT  55.81 52.31 56.14 52.05 ;
      RECT  54.89 62.23 58.89 62.68 ;
      RECT  54.89 56.94 58.89 57.35 ;
      RECT  55.77 58.06 56.1 58.21 ;
      RECT  57.79 57.35 58.09 57.76 ;
      RECT  55.79 58.21 56.08 58.37 ;
      RECT  55.74 57.35 56.03 57.82 ;
      RECT  56.45 57.58 56.77 57.9 ;
      RECT  57.63 61.97 57.95 62.23 ;
      RECT  56.51 60.18 56.8 60.47 ;
      RECT  56.96 57.58 57.28 57.9 ;
      RECT  56.93 60.72 57.22 61.01 ;
      RECT  55.81 61.97 56.14 62.23 ;
      RECT  54.89 62.69 58.89 62.24 ;
      RECT  54.89 67.98 58.89 67.57 ;
      RECT  55.77 66.86 56.1 66.71 ;
      RECT  57.79 67.57 58.09 67.16 ;
      RECT  55.79 66.71 56.08 66.55 ;
      RECT  55.74 67.57 56.03 67.1 ;
      RECT  56.45 67.34 56.77 67.02 ;
      RECT  57.63 62.95 57.95 62.69 ;
      RECT  56.51 64.74 56.8 64.45 ;
      RECT  56.96 67.34 57.28 67.02 ;
      RECT  56.93 64.2 57.22 63.91 ;
      RECT  55.81 62.95 56.14 62.69 ;
      RECT  54.89 72.87 58.89 73.32 ;
      RECT  54.89 67.58 58.89 67.99 ;
      RECT  55.77 68.7 56.1 68.85 ;
      RECT  57.79 67.99 58.09 68.4 ;
      RECT  55.79 68.85 56.08 69.01 ;
      RECT  55.74 67.99 56.03 68.46 ;
      RECT  56.45 68.22 56.77 68.54 ;
      RECT  57.63 72.61 57.95 72.87 ;
      RECT  56.51 70.82 56.8 71.11 ;
      RECT  56.96 68.22 57.28 68.54 ;
      RECT  56.93 71.36 57.22 71.65 ;
      RECT  55.81 72.61 56.14 72.87 ;
      RECT  54.89 73.33 58.89 72.88 ;
      RECT  54.89 78.62 58.89 78.21 ;
      RECT  55.77 77.5 56.1 77.35 ;
      RECT  57.79 78.21 58.09 77.8 ;
      RECT  55.79 77.35 56.08 77.19 ;
      RECT  55.74 78.21 56.03 77.74 ;
      RECT  56.45 77.98 56.77 77.66 ;
      RECT  57.63 73.59 57.95 73.33 ;
      RECT  56.51 75.38 56.8 75.09 ;
      RECT  56.96 77.98 57.28 77.66 ;
      RECT  56.93 74.84 57.22 74.55 ;
      RECT  55.81 73.59 56.14 73.33 ;
      RECT  54.89 83.51 58.89 83.96 ;
      RECT  54.89 78.22 58.89 78.63 ;
      RECT  55.77 79.34 56.1 79.49 ;
      RECT  57.79 78.63 58.09 79.04 ;
      RECT  55.79 79.49 56.08 79.65 ;
      RECT  55.74 78.63 56.03 79.1 ;
      RECT  56.45 78.86 56.77 79.18 ;
      RECT  57.63 83.25 57.95 83.51 ;
      RECT  56.51 81.46 56.8 81.75 ;
      RECT  56.96 78.86 57.28 79.18 ;
      RECT  56.93 82.0 57.22 82.29 ;
      RECT  55.81 83.25 56.14 83.51 ;
      RECT  54.89 83.97 58.89 83.52 ;
      RECT  54.89 89.26 58.89 88.85 ;
      RECT  55.77 88.14 56.1 87.99 ;
      RECT  57.79 88.85 58.09 88.44 ;
      RECT  55.79 87.99 56.08 87.83 ;
      RECT  55.74 88.85 56.03 88.38 ;
      RECT  56.45 88.62 56.77 88.3 ;
      RECT  57.63 84.23 57.95 83.97 ;
      RECT  56.51 86.02 56.8 85.73 ;
      RECT  56.96 88.62 57.28 88.3 ;
      RECT  56.93 85.48 57.22 85.19 ;
      RECT  55.81 84.23 56.14 83.97 ;
      RECT  54.89 94.15 58.89 94.6 ;
      RECT  54.89 88.86 58.89 89.27 ;
      RECT  55.77 89.98 56.1 90.13 ;
      RECT  57.79 89.27 58.09 89.68 ;
      RECT  55.79 90.13 56.08 90.29 ;
      RECT  55.74 89.27 56.03 89.74 ;
      RECT  56.45 89.5 56.77 89.82 ;
      RECT  57.63 93.89 57.95 94.15 ;
      RECT  56.51 92.1 56.8 92.39 ;
      RECT  56.96 89.5 57.28 89.82 ;
      RECT  56.93 92.64 57.22 92.93 ;
      RECT  55.81 93.89 56.14 94.15 ;
      RECT  54.89 94.61 58.89 94.16 ;
      RECT  54.89 99.9 58.89 99.49 ;
      RECT  55.77 98.78 56.1 98.63 ;
      RECT  57.79 99.49 58.09 99.08 ;
      RECT  55.79 98.63 56.08 98.47 ;
      RECT  55.74 99.49 56.03 99.02 ;
      RECT  56.45 99.26 56.77 98.94 ;
      RECT  57.63 94.87 57.95 94.61 ;
      RECT  56.51 96.66 56.8 96.37 ;
      RECT  56.96 99.26 57.28 98.94 ;
      RECT  56.93 96.12 57.22 95.83 ;
      RECT  55.81 94.87 56.14 94.61 ;
      RECT  54.89 104.79 58.89 105.24 ;
      RECT  54.89 99.5 58.89 99.91 ;
      RECT  55.77 100.62 56.1 100.77 ;
      RECT  57.79 99.91 58.09 100.32 ;
      RECT  55.79 100.77 56.08 100.93 ;
      RECT  55.74 99.91 56.03 100.38 ;
      RECT  56.45 100.14 56.77 100.46 ;
      RECT  57.63 104.53 57.95 104.79 ;
      RECT  56.51 102.74 56.8 103.03 ;
      RECT  56.96 100.14 57.28 100.46 ;
      RECT  56.93 103.28 57.22 103.57 ;
      RECT  55.81 104.53 56.14 104.79 ;
      RECT  54.89 105.25 58.89 104.8 ;
      RECT  54.89 110.54 58.89 110.13 ;
      RECT  55.77 109.42 56.1 109.27 ;
      RECT  57.79 110.13 58.09 109.72 ;
      RECT  55.79 109.27 56.08 109.11 ;
      RECT  55.74 110.13 56.03 109.66 ;
      RECT  56.45 109.9 56.77 109.58 ;
      RECT  57.63 105.51 57.95 105.25 ;
      RECT  56.51 107.3 56.8 107.01 ;
      RECT  56.96 109.9 57.28 109.58 ;
      RECT  56.93 106.76 57.22 106.47 ;
      RECT  55.81 105.51 56.14 105.25 ;
      RECT  54.89 115.43 58.89 115.88 ;
      RECT  54.89 110.14 58.89 110.55 ;
      RECT  55.77 111.26 56.1 111.41 ;
      RECT  57.79 110.55 58.09 110.96 ;
      RECT  55.79 111.41 56.08 111.57 ;
      RECT  55.74 110.55 56.03 111.02 ;
      RECT  56.45 110.78 56.77 111.1 ;
      RECT  57.63 115.17 57.95 115.43 ;
      RECT  56.51 113.38 56.8 113.67 ;
      RECT  56.96 110.78 57.28 111.1 ;
      RECT  56.93 113.92 57.22 114.21 ;
      RECT  55.81 115.17 56.14 115.43 ;
      RECT  54.89 115.89 58.89 115.44 ;
      RECT  54.89 121.18 58.89 120.77 ;
      RECT  55.77 120.06 56.1 119.91 ;
      RECT  57.79 120.77 58.09 120.36 ;
      RECT  55.79 119.91 56.08 119.75 ;
      RECT  55.74 120.77 56.03 120.3 ;
      RECT  56.45 120.54 56.77 120.22 ;
      RECT  57.63 116.15 57.95 115.89 ;
      RECT  56.51 117.94 56.8 117.65 ;
      RECT  56.96 120.54 57.28 120.22 ;
      RECT  56.93 117.4 57.22 117.11 ;
      RECT  55.81 116.15 56.14 115.89 ;
      RECT  58.89 40.95 62.89 41.4 ;
      RECT  58.89 35.66 62.89 36.07 ;
      RECT  59.77 36.78 60.1 36.93 ;
      RECT  61.79 36.07 62.09 36.48 ;
      RECT  59.79 36.93 60.08 37.09 ;
      RECT  59.74 36.07 60.03 36.54 ;
      RECT  60.45 36.3 60.77 36.62 ;
      RECT  61.63 40.69 61.95 40.95 ;
      RECT  60.51 38.9 60.8 39.19 ;
      RECT  60.96 36.3 61.28 36.62 ;
      RECT  60.93 39.44 61.22 39.73 ;
      RECT  59.81 40.69 60.14 40.95 ;
      RECT  58.89 41.41 62.89 40.96 ;
      RECT  58.89 46.7 62.89 46.29 ;
      RECT  59.77 45.58 60.1 45.43 ;
      RECT  61.79 46.29 62.09 45.88 ;
      RECT  59.79 45.43 60.08 45.27 ;
      RECT  59.74 46.29 60.03 45.82 ;
      RECT  60.45 46.06 60.77 45.74 ;
      RECT  61.63 41.67 61.95 41.41 ;
      RECT  60.51 43.46 60.8 43.17 ;
      RECT  60.96 46.06 61.28 45.74 ;
      RECT  60.93 42.92 61.22 42.63 ;
      RECT  59.81 41.67 60.14 41.41 ;
      RECT  58.89 51.59 62.89 52.04 ;
      RECT  58.89 46.3 62.89 46.71 ;
      RECT  59.77 47.42 60.1 47.57 ;
      RECT  61.79 46.71 62.09 47.12 ;
      RECT  59.79 47.57 60.08 47.73 ;
      RECT  59.74 46.71 60.03 47.18 ;
      RECT  60.45 46.94 60.77 47.26 ;
      RECT  61.63 51.33 61.95 51.59 ;
      RECT  60.51 49.54 60.8 49.83 ;
      RECT  60.96 46.94 61.28 47.26 ;
      RECT  60.93 50.08 61.22 50.37 ;
      RECT  59.81 51.33 60.14 51.59 ;
      RECT  58.89 52.05 62.89 51.6 ;
      RECT  58.89 57.34 62.89 56.93 ;
      RECT  59.77 56.22 60.1 56.07 ;
      RECT  61.79 56.93 62.09 56.52 ;
      RECT  59.79 56.07 60.08 55.91 ;
      RECT  59.74 56.93 60.03 56.46 ;
      RECT  60.45 56.7 60.77 56.38 ;
      RECT  61.63 52.31 61.95 52.05 ;
      RECT  60.51 54.1 60.8 53.81 ;
      RECT  60.96 56.7 61.28 56.38 ;
      RECT  60.93 53.56 61.22 53.27 ;
      RECT  59.81 52.31 60.14 52.05 ;
      RECT  58.89 62.23 62.89 62.68 ;
      RECT  58.89 56.94 62.89 57.35 ;
      RECT  59.77 58.06 60.1 58.21 ;
      RECT  61.79 57.35 62.09 57.76 ;
      RECT  59.79 58.21 60.08 58.37 ;
      RECT  59.74 57.35 60.03 57.82 ;
      RECT  60.45 57.58 60.77 57.9 ;
      RECT  61.63 61.97 61.95 62.23 ;
      RECT  60.51 60.18 60.8 60.47 ;
      RECT  60.96 57.58 61.28 57.9 ;
      RECT  60.93 60.72 61.22 61.01 ;
      RECT  59.81 61.97 60.14 62.23 ;
      RECT  58.89 62.69 62.89 62.24 ;
      RECT  58.89 67.98 62.89 67.57 ;
      RECT  59.77 66.86 60.1 66.71 ;
      RECT  61.79 67.57 62.09 67.16 ;
      RECT  59.79 66.71 60.08 66.55 ;
      RECT  59.74 67.57 60.03 67.1 ;
      RECT  60.45 67.34 60.77 67.02 ;
      RECT  61.63 62.95 61.95 62.69 ;
      RECT  60.51 64.74 60.8 64.45 ;
      RECT  60.96 67.34 61.28 67.02 ;
      RECT  60.93 64.2 61.22 63.91 ;
      RECT  59.81 62.95 60.14 62.69 ;
      RECT  58.89 72.87 62.89 73.32 ;
      RECT  58.89 67.58 62.89 67.99 ;
      RECT  59.77 68.7 60.1 68.85 ;
      RECT  61.79 67.99 62.09 68.4 ;
      RECT  59.79 68.85 60.08 69.01 ;
      RECT  59.74 67.99 60.03 68.46 ;
      RECT  60.45 68.22 60.77 68.54 ;
      RECT  61.63 72.61 61.95 72.87 ;
      RECT  60.51 70.82 60.8 71.11 ;
      RECT  60.96 68.22 61.28 68.54 ;
      RECT  60.93 71.36 61.22 71.65 ;
      RECT  59.81 72.61 60.14 72.87 ;
      RECT  58.89 73.33 62.89 72.88 ;
      RECT  58.89 78.62 62.89 78.21 ;
      RECT  59.77 77.5 60.1 77.35 ;
      RECT  61.79 78.21 62.09 77.8 ;
      RECT  59.79 77.35 60.08 77.19 ;
      RECT  59.74 78.21 60.03 77.74 ;
      RECT  60.45 77.98 60.77 77.66 ;
      RECT  61.63 73.59 61.95 73.33 ;
      RECT  60.51 75.38 60.8 75.09 ;
      RECT  60.96 77.98 61.28 77.66 ;
      RECT  60.93 74.84 61.22 74.55 ;
      RECT  59.81 73.59 60.14 73.33 ;
      RECT  58.89 83.51 62.89 83.96 ;
      RECT  58.89 78.22 62.89 78.63 ;
      RECT  59.77 79.34 60.1 79.49 ;
      RECT  61.79 78.63 62.09 79.04 ;
      RECT  59.79 79.49 60.08 79.65 ;
      RECT  59.74 78.63 60.03 79.1 ;
      RECT  60.45 78.86 60.77 79.18 ;
      RECT  61.63 83.25 61.95 83.51 ;
      RECT  60.51 81.46 60.8 81.75 ;
      RECT  60.96 78.86 61.28 79.18 ;
      RECT  60.93 82.0 61.22 82.29 ;
      RECT  59.81 83.25 60.14 83.51 ;
      RECT  58.89 83.97 62.89 83.52 ;
      RECT  58.89 89.26 62.89 88.85 ;
      RECT  59.77 88.14 60.1 87.99 ;
      RECT  61.79 88.85 62.09 88.44 ;
      RECT  59.79 87.99 60.08 87.83 ;
      RECT  59.74 88.85 60.03 88.38 ;
      RECT  60.45 88.62 60.77 88.3 ;
      RECT  61.63 84.23 61.95 83.97 ;
      RECT  60.51 86.02 60.8 85.73 ;
      RECT  60.96 88.62 61.28 88.3 ;
      RECT  60.93 85.48 61.22 85.19 ;
      RECT  59.81 84.23 60.14 83.97 ;
      RECT  58.89 94.15 62.89 94.6 ;
      RECT  58.89 88.86 62.89 89.27 ;
      RECT  59.77 89.98 60.1 90.13 ;
      RECT  61.79 89.27 62.09 89.68 ;
      RECT  59.79 90.13 60.08 90.29 ;
      RECT  59.74 89.27 60.03 89.74 ;
      RECT  60.45 89.5 60.77 89.82 ;
      RECT  61.63 93.89 61.95 94.15 ;
      RECT  60.51 92.1 60.8 92.39 ;
      RECT  60.96 89.5 61.28 89.82 ;
      RECT  60.93 92.64 61.22 92.93 ;
      RECT  59.81 93.89 60.14 94.15 ;
      RECT  58.89 94.61 62.89 94.16 ;
      RECT  58.89 99.9 62.89 99.49 ;
      RECT  59.77 98.78 60.1 98.63 ;
      RECT  61.79 99.49 62.09 99.08 ;
      RECT  59.79 98.63 60.08 98.47 ;
      RECT  59.74 99.49 60.03 99.02 ;
      RECT  60.45 99.26 60.77 98.94 ;
      RECT  61.63 94.87 61.95 94.61 ;
      RECT  60.51 96.66 60.8 96.37 ;
      RECT  60.96 99.26 61.28 98.94 ;
      RECT  60.93 96.12 61.22 95.83 ;
      RECT  59.81 94.87 60.14 94.61 ;
      RECT  58.89 104.79 62.89 105.24 ;
      RECT  58.89 99.5 62.89 99.91 ;
      RECT  59.77 100.62 60.1 100.77 ;
      RECT  61.79 99.91 62.09 100.32 ;
      RECT  59.79 100.77 60.08 100.93 ;
      RECT  59.74 99.91 60.03 100.38 ;
      RECT  60.45 100.14 60.77 100.46 ;
      RECT  61.63 104.53 61.95 104.79 ;
      RECT  60.51 102.74 60.8 103.03 ;
      RECT  60.96 100.14 61.28 100.46 ;
      RECT  60.93 103.28 61.22 103.57 ;
      RECT  59.81 104.53 60.14 104.79 ;
      RECT  58.89 105.25 62.89 104.8 ;
      RECT  58.89 110.54 62.89 110.13 ;
      RECT  59.77 109.42 60.1 109.27 ;
      RECT  61.79 110.13 62.09 109.72 ;
      RECT  59.79 109.27 60.08 109.11 ;
      RECT  59.74 110.13 60.03 109.66 ;
      RECT  60.45 109.9 60.77 109.58 ;
      RECT  61.63 105.51 61.95 105.25 ;
      RECT  60.51 107.3 60.8 107.01 ;
      RECT  60.96 109.9 61.28 109.58 ;
      RECT  60.93 106.76 61.22 106.47 ;
      RECT  59.81 105.51 60.14 105.25 ;
      RECT  58.89 115.43 62.89 115.88 ;
      RECT  58.89 110.14 62.89 110.55 ;
      RECT  59.77 111.26 60.1 111.41 ;
      RECT  61.79 110.55 62.09 110.96 ;
      RECT  59.79 111.41 60.08 111.57 ;
      RECT  59.74 110.55 60.03 111.02 ;
      RECT  60.45 110.78 60.77 111.1 ;
      RECT  61.63 115.17 61.95 115.43 ;
      RECT  60.51 113.38 60.8 113.67 ;
      RECT  60.96 110.78 61.28 111.1 ;
      RECT  60.93 113.92 61.22 114.21 ;
      RECT  59.81 115.17 60.14 115.43 ;
      RECT  58.89 115.89 62.89 115.44 ;
      RECT  58.89 121.18 62.89 120.77 ;
      RECT  59.77 120.06 60.1 119.91 ;
      RECT  61.79 120.77 62.09 120.36 ;
      RECT  59.79 119.91 60.08 119.75 ;
      RECT  59.74 120.77 60.03 120.3 ;
      RECT  60.45 120.54 60.77 120.22 ;
      RECT  61.63 116.15 61.95 115.89 ;
      RECT  60.51 117.94 60.8 117.65 ;
      RECT  60.96 120.54 61.28 120.22 ;
      RECT  60.93 117.4 61.22 117.11 ;
      RECT  59.81 116.15 60.14 115.89 ;
      RECT  54.89 36.93 62.89 37.09 ;
      RECT  54.89 45.27 62.89 45.43 ;
      RECT  54.89 47.57 62.89 47.73 ;
      RECT  54.89 55.91 62.89 56.07 ;
      RECT  54.89 58.21 62.89 58.37 ;
      RECT  54.89 66.55 62.89 66.71 ;
      RECT  54.89 68.85 62.89 69.01 ;
      RECT  54.89 77.19 62.89 77.35 ;
      RECT  54.89 79.49 62.89 79.65 ;
      RECT  54.89 87.83 62.89 87.99 ;
      RECT  54.89 90.13 62.89 90.29 ;
      RECT  54.89 98.47 62.89 98.63 ;
      RECT  54.89 100.77 62.89 100.93 ;
      RECT  54.89 109.11 62.89 109.27 ;
      RECT  54.89 111.41 62.89 111.57 ;
      RECT  54.89 119.75 62.89 119.91 ;
      RECT  54.89 40.96 58.89 41.41 ;
      RECT  54.89 40.95 58.89 41.4 ;
      RECT  54.89 104.8 58.89 105.25 ;
      RECT  58.89 104.79 62.89 105.24 ;
      RECT  54.89 72.88 58.89 73.33 ;
      RECT  54.89 94.16 58.89 94.61 ;
      RECT  58.89 72.87 62.89 73.32 ;
      RECT  54.89 83.52 58.89 83.97 ;
      RECT  58.89 72.88 62.89 73.33 ;
      RECT  54.89 62.23 58.89 62.68 ;
      RECT  58.89 115.43 62.89 115.88 ;
      RECT  54.89 94.15 58.89 94.6 ;
      RECT  58.89 62.24 62.89 62.69 ;
      RECT  58.89 51.59 62.89 52.04 ;
      RECT  58.89 40.95 62.89 41.4 ;
      RECT  54.89 104.79 58.89 105.24 ;
      RECT  54.89 51.6 58.89 52.05 ;
      RECT  58.89 94.15 62.89 94.6 ;
      RECT  58.89 40.96 62.89 41.41 ;
      RECT  58.89 104.8 62.89 105.25 ;
      RECT  58.89 62.23 62.89 62.68 ;
      RECT  58.89 51.6 62.89 52.05 ;
      RECT  54.89 62.24 58.89 62.69 ;
      RECT  58.89 83.52 62.89 83.97 ;
      RECT  54.89 72.87 58.89 73.32 ;
      RECT  58.89 83.51 62.89 83.96 ;
      RECT  54.89 83.51 58.89 83.96 ;
      RECT  58.89 94.16 62.89 94.61 ;
      RECT  54.89 115.43 58.89 115.88 ;
      RECT  54.89 51.59 58.89 52.04 ;
      RECT  58.89 115.44 62.89 115.89 ;
      RECT  54.89 115.44 58.89 115.89 ;
      RECT  54.89 110.13 58.89 110.54 ;
      RECT  58.89 67.57 62.89 67.98 ;
      RECT  54.89 120.77 58.89 121.18 ;
      RECT  54.89 67.57 58.89 67.98 ;
      RECT  58.89 78.21 62.89 78.62 ;
      RECT  58.89 46.3 62.89 46.71 ;
      RECT  54.89 110.14 58.89 110.55 ;
      RECT  58.89 56.93 62.89 57.34 ;
      RECT  58.89 67.58 62.89 67.99 ;
      RECT  58.89 120.77 62.89 121.18 ;
      RECT  54.89 56.94 58.89 57.35 ;
      RECT  54.89 88.86 58.89 89.27 ;
      RECT  54.89 56.93 58.89 57.34 ;
      RECT  58.89 88.86 62.89 89.27 ;
      RECT  58.89 110.13 62.89 110.54 ;
      RECT  54.89 88.85 58.89 89.26 ;
      RECT  58.89 88.85 62.89 89.26 ;
      RECT  58.89 99.5 62.89 99.91 ;
      RECT  58.89 78.22 62.89 78.63 ;
      RECT  54.89 35.66 58.89 36.07 ;
      RECT  54.89 99.5 58.89 99.91 ;
      RECT  58.89 35.66 62.89 36.07 ;
      RECT  54.89 78.22 58.89 78.63 ;
      RECT  54.89 67.58 58.89 67.99 ;
      RECT  54.89 78.21 58.89 78.62 ;
      RECT  54.89 46.3 58.89 46.71 ;
      RECT  58.89 99.49 62.89 99.9 ;
      RECT  54.89 99.49 58.89 99.9 ;
      RECT  58.89 56.94 62.89 57.35 ;
      RECT  54.89 46.29 58.89 46.7 ;
      RECT  58.89 46.29 62.89 46.7 ;
      RECT  58.89 110.14 62.89 110.55 ;
      RECT  50.89 30.31 54.89 30.76 ;
      RECT  50.89 25.02 54.89 25.43 ;
      RECT  51.77 26.14 52.1 26.29 ;
      RECT  53.79 25.43 54.09 25.84 ;
      RECT  51.79 26.29 52.08 26.45 ;
      RECT  51.74 25.43 52.03 25.9 ;
      RECT  53.63 30.05 53.95 30.31 ;
      RECT  52.51 28.26 52.8 28.55 ;
      RECT  52.93 28.8 53.22 29.09 ;
      RECT  51.81 30.05 52.14 30.31 ;
      RECT  50.89 30.77 54.89 30.32 ;
      RECT  50.89 36.06 54.89 35.65 ;
      RECT  51.77 34.94 52.1 34.79 ;
      RECT  53.79 35.65 54.09 35.24 ;
      RECT  51.79 34.79 52.08 34.63 ;
      RECT  51.74 35.65 52.03 35.18 ;
      RECT  52.45 35.42 52.77 35.1 ;
      RECT  53.63 31.03 53.95 30.77 ;
      RECT  52.51 32.82 52.8 32.53 ;
      RECT  52.96 35.42 53.28 35.1 ;
      RECT  53.02 31.02 53.34 30.77 ;
      RECT  52.93 32.28 53.22 31.99 ;
      RECT  51.81 31.03 52.14 30.77 ;
      RECT  50.89 40.95 54.89 41.4 ;
      RECT  50.89 35.66 54.89 36.07 ;
      RECT  51.77 36.78 52.1 36.93 ;
      RECT  53.79 36.07 54.09 36.48 ;
      RECT  51.79 36.93 52.08 37.09 ;
      RECT  51.74 36.07 52.03 36.54 ;
      RECT  52.45 36.3 52.77 36.62 ;
      RECT  53.63 40.69 53.95 40.95 ;
      RECT  52.51 38.9 52.8 39.19 ;
      RECT  52.96 36.3 53.28 36.62 ;
      RECT  53.02 40.7 53.34 40.95 ;
      RECT  52.93 39.44 53.22 39.73 ;
      RECT  51.81 40.69 52.14 40.95 ;
      RECT  50.89 41.41 54.89 40.96 ;
      RECT  50.89 46.7 54.89 46.29 ;
      RECT  51.77 45.58 52.1 45.43 ;
      RECT  53.79 46.29 54.09 45.88 ;
      RECT  51.79 45.43 52.08 45.27 ;
      RECT  51.74 46.29 52.03 45.82 ;
      RECT  52.45 46.06 52.77 45.74 ;
      RECT  53.63 41.67 53.95 41.41 ;
      RECT  52.51 43.46 52.8 43.17 ;
      RECT  52.96 46.06 53.28 45.74 ;
      RECT  53.02 41.66 53.34 41.41 ;
      RECT  52.93 42.92 53.22 42.63 ;
      RECT  51.81 41.67 52.14 41.41 ;
      RECT  50.89 51.59 54.89 52.04 ;
      RECT  50.89 46.3 54.89 46.71 ;
      RECT  51.77 47.42 52.1 47.57 ;
      RECT  53.79 46.71 54.09 47.12 ;
      RECT  51.79 47.57 52.08 47.73 ;
      RECT  51.74 46.71 52.03 47.18 ;
      RECT  52.45 46.94 52.77 47.26 ;
      RECT  53.63 51.33 53.95 51.59 ;
      RECT  52.51 49.54 52.8 49.83 ;
      RECT  52.96 46.94 53.28 47.26 ;
      RECT  53.02 51.34 53.34 51.59 ;
      RECT  52.93 50.08 53.22 50.37 ;
      RECT  51.81 51.33 52.14 51.59 ;
      RECT  50.89 52.05 54.89 51.6 ;
      RECT  50.89 57.34 54.89 56.93 ;
      RECT  51.77 56.22 52.1 56.07 ;
      RECT  53.79 56.93 54.09 56.52 ;
      RECT  51.79 56.07 52.08 55.91 ;
      RECT  51.74 56.93 52.03 56.46 ;
      RECT  52.45 56.7 52.77 56.38 ;
      RECT  53.63 52.31 53.95 52.05 ;
      RECT  52.51 54.1 52.8 53.81 ;
      RECT  52.96 56.7 53.28 56.38 ;
      RECT  53.02 52.3 53.34 52.05 ;
      RECT  52.93 53.56 53.22 53.27 ;
      RECT  51.81 52.31 52.14 52.05 ;
      RECT  50.89 62.23 54.89 62.68 ;
      RECT  50.89 56.94 54.89 57.35 ;
      RECT  51.77 58.06 52.1 58.21 ;
      RECT  53.79 57.35 54.09 57.76 ;
      RECT  51.79 58.21 52.08 58.37 ;
      RECT  51.74 57.35 52.03 57.82 ;
      RECT  52.45 57.58 52.77 57.9 ;
      RECT  53.63 61.97 53.95 62.23 ;
      RECT  52.51 60.18 52.8 60.47 ;
      RECT  52.96 57.58 53.28 57.9 ;
      RECT  53.02 61.98 53.34 62.23 ;
      RECT  52.93 60.72 53.22 61.01 ;
      RECT  51.81 61.97 52.14 62.23 ;
      RECT  50.89 62.69 54.89 62.24 ;
      RECT  50.89 67.98 54.89 67.57 ;
      RECT  51.77 66.86 52.1 66.71 ;
      RECT  53.79 67.57 54.09 67.16 ;
      RECT  51.79 66.71 52.08 66.55 ;
      RECT  51.74 67.57 52.03 67.1 ;
      RECT  52.45 67.34 52.77 67.02 ;
      RECT  53.63 62.95 53.95 62.69 ;
      RECT  52.51 64.74 52.8 64.45 ;
      RECT  52.96 67.34 53.28 67.02 ;
      RECT  53.02 62.94 53.34 62.69 ;
      RECT  52.93 64.2 53.22 63.91 ;
      RECT  51.81 62.95 52.14 62.69 ;
      RECT  50.89 72.87 54.89 73.32 ;
      RECT  50.89 67.58 54.89 67.99 ;
      RECT  51.77 68.7 52.1 68.85 ;
      RECT  53.79 67.99 54.09 68.4 ;
      RECT  51.79 68.85 52.08 69.01 ;
      RECT  51.74 67.99 52.03 68.46 ;
      RECT  52.45 68.22 52.77 68.54 ;
      RECT  53.63 72.61 53.95 72.87 ;
      RECT  52.51 70.82 52.8 71.11 ;
      RECT  52.96 68.22 53.28 68.54 ;
      RECT  53.02 72.62 53.34 72.87 ;
      RECT  52.93 71.36 53.22 71.65 ;
      RECT  51.81 72.61 52.14 72.87 ;
      RECT  50.89 73.33 54.89 72.88 ;
      RECT  50.89 78.62 54.89 78.21 ;
      RECT  51.77 77.5 52.1 77.35 ;
      RECT  53.79 78.21 54.09 77.8 ;
      RECT  51.79 77.35 52.08 77.19 ;
      RECT  51.74 78.21 52.03 77.74 ;
      RECT  52.45 77.98 52.77 77.66 ;
      RECT  53.63 73.59 53.95 73.33 ;
      RECT  52.51 75.38 52.8 75.09 ;
      RECT  52.96 77.98 53.28 77.66 ;
      RECT  53.02 73.58 53.34 73.33 ;
      RECT  52.93 74.84 53.22 74.55 ;
      RECT  51.81 73.59 52.14 73.33 ;
      RECT  50.89 83.51 54.89 83.96 ;
      RECT  50.89 78.22 54.89 78.63 ;
      RECT  51.77 79.34 52.1 79.49 ;
      RECT  53.79 78.63 54.09 79.04 ;
      RECT  51.79 79.49 52.08 79.65 ;
      RECT  51.74 78.63 52.03 79.1 ;
      RECT  52.45 78.86 52.77 79.18 ;
      RECT  53.63 83.25 53.95 83.51 ;
      RECT  52.51 81.46 52.8 81.75 ;
      RECT  52.96 78.86 53.28 79.18 ;
      RECT  53.02 83.26 53.34 83.51 ;
      RECT  52.93 82.0 53.22 82.29 ;
      RECT  51.81 83.25 52.14 83.51 ;
      RECT  50.89 83.97 54.89 83.52 ;
      RECT  50.89 89.26 54.89 88.85 ;
      RECT  51.77 88.14 52.1 87.99 ;
      RECT  53.79 88.85 54.09 88.44 ;
      RECT  51.79 87.99 52.08 87.83 ;
      RECT  51.74 88.85 52.03 88.38 ;
      RECT  52.45 88.62 52.77 88.3 ;
      RECT  53.63 84.23 53.95 83.97 ;
      RECT  52.51 86.02 52.8 85.73 ;
      RECT  52.96 88.62 53.28 88.3 ;
      RECT  53.02 84.22 53.34 83.97 ;
      RECT  52.93 85.48 53.22 85.19 ;
      RECT  51.81 84.23 52.14 83.97 ;
      RECT  50.89 94.15 54.89 94.6 ;
      RECT  50.89 88.86 54.89 89.27 ;
      RECT  51.77 89.98 52.1 90.13 ;
      RECT  53.79 89.27 54.09 89.68 ;
      RECT  51.79 90.13 52.08 90.29 ;
      RECT  51.74 89.27 52.03 89.74 ;
      RECT  52.45 89.5 52.77 89.82 ;
      RECT  53.63 93.89 53.95 94.15 ;
      RECT  52.51 92.1 52.8 92.39 ;
      RECT  52.96 89.5 53.28 89.82 ;
      RECT  53.02 93.9 53.34 94.15 ;
      RECT  52.93 92.64 53.22 92.93 ;
      RECT  51.81 93.89 52.14 94.15 ;
      RECT  50.89 94.61 54.89 94.16 ;
      RECT  50.89 99.9 54.89 99.49 ;
      RECT  51.77 98.78 52.1 98.63 ;
      RECT  53.79 99.49 54.09 99.08 ;
      RECT  51.79 98.63 52.08 98.47 ;
      RECT  51.74 99.49 52.03 99.02 ;
      RECT  52.45 99.26 52.77 98.94 ;
      RECT  53.63 94.87 53.95 94.61 ;
      RECT  52.51 96.66 52.8 96.37 ;
      RECT  52.96 99.26 53.28 98.94 ;
      RECT  53.02 94.86 53.34 94.61 ;
      RECT  52.93 96.12 53.22 95.83 ;
      RECT  51.81 94.87 52.14 94.61 ;
      RECT  50.89 104.79 54.89 105.24 ;
      RECT  50.89 99.5 54.89 99.91 ;
      RECT  51.77 100.62 52.1 100.77 ;
      RECT  53.79 99.91 54.09 100.32 ;
      RECT  51.79 100.77 52.08 100.93 ;
      RECT  51.74 99.91 52.03 100.38 ;
      RECT  52.45 100.14 52.77 100.46 ;
      RECT  53.63 104.53 53.95 104.79 ;
      RECT  52.51 102.74 52.8 103.03 ;
      RECT  52.96 100.14 53.28 100.46 ;
      RECT  53.02 104.54 53.34 104.79 ;
      RECT  52.93 103.28 53.22 103.57 ;
      RECT  51.81 104.53 52.14 104.79 ;
      RECT  50.89 105.25 54.89 104.8 ;
      RECT  50.89 110.54 54.89 110.13 ;
      RECT  51.77 109.42 52.1 109.27 ;
      RECT  53.79 110.13 54.09 109.72 ;
      RECT  51.79 109.27 52.08 109.11 ;
      RECT  51.74 110.13 52.03 109.66 ;
      RECT  52.45 109.9 52.77 109.58 ;
      RECT  53.63 105.51 53.95 105.25 ;
      RECT  52.51 107.3 52.8 107.01 ;
      RECT  52.96 109.9 53.28 109.58 ;
      RECT  53.02 105.5 53.34 105.25 ;
      RECT  52.93 106.76 53.22 106.47 ;
      RECT  51.81 105.51 52.14 105.25 ;
      RECT  50.89 115.43 54.89 115.88 ;
      RECT  50.89 110.14 54.89 110.55 ;
      RECT  51.77 111.26 52.1 111.41 ;
      RECT  53.79 110.55 54.09 110.96 ;
      RECT  51.79 111.41 52.08 111.57 ;
      RECT  51.74 110.55 52.03 111.02 ;
      RECT  52.45 110.78 52.77 111.1 ;
      RECT  53.63 115.17 53.95 115.43 ;
      RECT  52.51 113.38 52.8 113.67 ;
      RECT  52.96 110.78 53.28 111.1 ;
      RECT  53.02 115.18 53.34 115.43 ;
      RECT  52.93 113.92 53.22 114.21 ;
      RECT  51.81 115.17 52.14 115.43 ;
      RECT  50.89 115.89 54.89 115.44 ;
      RECT  50.89 121.18 54.89 120.77 ;
      RECT  51.77 120.06 52.1 119.91 ;
      RECT  53.79 120.77 54.09 120.36 ;
      RECT  51.79 119.91 52.08 119.75 ;
      RECT  51.74 120.77 52.03 120.3 ;
      RECT  52.45 120.54 52.77 120.22 ;
      RECT  53.63 116.15 53.95 115.89 ;
      RECT  52.51 117.94 52.8 117.65 ;
      RECT  52.96 120.54 53.28 120.22 ;
      RECT  53.02 116.14 53.34 115.89 ;
      RECT  52.93 117.4 53.22 117.11 ;
      RECT  51.81 116.15 52.14 115.89 ;
      RECT  50.89 126.07 54.89 126.52 ;
      RECT  50.89 120.78 54.89 121.19 ;
      RECT  51.77 121.9 52.1 122.05 ;
      RECT  53.79 121.19 54.09 121.6 ;
      RECT  51.79 122.05 52.08 122.21 ;
      RECT  51.74 121.19 52.03 121.66 ;
      RECT  53.63 125.81 53.95 126.07 ;
      RECT  52.51 124.02 52.8 124.31 ;
      RECT  52.93 124.56 53.22 124.85 ;
      RECT  51.81 125.81 52.14 126.07 ;
      RECT  50.89 26.29 54.89 26.45 ;
      RECT  50.89 34.63 54.89 34.79 ;
      RECT  50.89 36.93 54.89 37.09 ;
      RECT  50.89 45.27 54.89 45.43 ;
      RECT  50.89 47.57 54.89 47.73 ;
      RECT  50.89 55.91 54.89 56.07 ;
      RECT  50.89 58.21 54.89 58.37 ;
      RECT  50.89 66.55 54.89 66.71 ;
      RECT  50.89 68.85 54.89 69.01 ;
      RECT  50.89 77.19 54.89 77.35 ;
      RECT  50.89 79.49 54.89 79.65 ;
      RECT  50.89 87.83 54.89 87.99 ;
      RECT  50.89 90.13 54.89 90.29 ;
      RECT  50.89 98.47 54.89 98.63 ;
      RECT  50.89 100.77 54.89 100.93 ;
      RECT  50.89 109.11 54.89 109.27 ;
      RECT  50.89 111.41 54.89 111.57 ;
      RECT  50.89 119.75 54.89 119.91 ;
      RECT  50.89 122.05 54.89 122.21 ;
      RECT  50.89 30.32 54.89 30.77 ;
      RECT  50.89 94.16 54.89 94.61 ;
      RECT  50.89 62.24 54.89 62.69 ;
      RECT  50.89 83.52 54.89 83.97 ;
      RECT  50.89 51.59 54.89 52.04 ;
      RECT  50.89 72.88 54.89 73.33 ;
      RECT  50.89 83.51 54.89 83.96 ;
      RECT  50.89 94.15 54.89 94.6 ;
      RECT  50.89 115.44 54.89 115.89 ;
      RECT  50.89 40.96 54.89 41.41 ;
      RECT  50.89 51.6 54.89 52.05 ;
      RECT  50.89 62.23 54.89 62.68 ;
      RECT  50.89 115.43 54.89 115.88 ;
      RECT  50.89 72.87 54.89 73.32 ;
      RECT  50.89 104.79 54.89 105.24 ;
      RECT  50.89 40.95 54.89 41.4 ;
      RECT  50.89 104.8 54.89 105.25 ;
      RECT  50.89 99.49 54.89 99.9 ;
      RECT  50.89 110.13 54.89 110.54 ;
      RECT  50.89 56.93 54.89 57.34 ;
      RECT  50.89 110.14 54.89 110.55 ;
      RECT  50.89 120.77 54.89 121.18 ;
      RECT  50.89 99.5 54.89 99.91 ;
      RECT  50.89 46.3 54.89 46.71 ;
      RECT  50.89 78.22 54.89 78.63 ;
      RECT  50.89 46.29 54.89 46.7 ;
      RECT  50.89 78.21 54.89 78.62 ;
      RECT  50.89 88.86 54.89 89.27 ;
      RECT  50.89 67.58 54.89 67.99 ;
      RECT  50.89 56.94 54.89 57.35 ;
      RECT  50.89 35.66 54.89 36.07 ;
      RECT  50.89 67.57 54.89 67.98 ;
      RECT  50.89 88.85 54.89 89.26 ;
      RECT  50.89 35.65 54.89 36.06 ;
      RECT  54.89 30.77 58.89 30.32 ;
      RECT  54.89 36.06 58.89 35.65 ;
      RECT  55.77 34.94 56.1 34.79 ;
      RECT  57.79 35.65 58.09 35.24 ;
      RECT  55.79 34.79 56.08 34.63 ;
      RECT  55.74 35.65 56.03 35.18 ;
      RECT  57.63 31.03 57.95 30.77 ;
      RECT  56.51 32.82 56.8 32.53 ;
      RECT  56.93 32.28 57.22 31.99 ;
      RECT  55.81 31.03 56.14 30.77 ;
      RECT  58.89 30.77 62.89 30.32 ;
      RECT  58.89 36.06 62.89 35.65 ;
      RECT  59.77 34.94 60.1 34.79 ;
      RECT  61.79 35.65 62.09 35.24 ;
      RECT  59.79 34.79 60.08 34.63 ;
      RECT  59.74 35.65 60.03 35.18 ;
      RECT  61.63 31.03 61.95 30.77 ;
      RECT  60.51 32.82 60.8 32.53 ;
      RECT  60.93 32.28 61.22 31.99 ;
      RECT  59.81 31.03 60.14 30.77 ;
      RECT  54.89 34.79 62.89 34.63 ;
      RECT  54.89 30.77 58.89 30.32 ;
      RECT  58.89 30.77 62.89 30.32 ;
      RECT  58.89 36.06 62.89 35.65 ;
      RECT  54.89 36.06 58.89 35.65 ;
      RECT  54.89 30.31 58.89 30.76 ;
      RECT  54.89 25.02 58.89 25.43 ;
      RECT  55.77 26.14 56.1 26.29 ;
      RECT  57.79 25.43 58.09 25.84 ;
      RECT  55.79 26.29 56.08 26.45 ;
      RECT  55.74 25.43 56.03 25.9 ;
      RECT  57.63 30.05 57.95 30.31 ;
      RECT  56.51 28.26 56.8 28.55 ;
      RECT  56.93 28.8 57.22 29.09 ;
      RECT  55.81 30.05 56.14 30.31 ;
      RECT  58.89 30.31 62.89 30.76 ;
      RECT  58.89 25.02 62.89 25.43 ;
      RECT  59.77 26.14 60.1 26.29 ;
      RECT  61.79 25.43 62.09 25.84 ;
      RECT  59.79 26.29 60.08 26.45 ;
      RECT  59.74 25.43 60.03 25.9 ;
      RECT  61.63 30.05 61.95 30.31 ;
      RECT  60.51 28.26 60.8 28.55 ;
      RECT  60.93 28.8 61.22 29.09 ;
      RECT  59.81 30.05 60.14 30.31 ;
      RECT  54.89 26.29 62.89 26.45 ;
      RECT  54.89 30.31 58.89 30.76 ;
      RECT  58.89 30.31 62.89 30.76 ;
      RECT  58.89 25.02 62.89 25.43 ;
      RECT  54.89 25.02 58.89 25.43 ;
      RECT  54.89 126.07 58.89 126.52 ;
      RECT  54.89 120.78 58.89 121.19 ;
      RECT  55.77 121.9 56.1 122.05 ;
      RECT  57.79 121.19 58.09 121.6 ;
      RECT  55.79 122.05 56.08 122.21 ;
      RECT  55.74 121.19 56.03 121.66 ;
      RECT  57.63 125.81 57.95 126.07 ;
      RECT  56.51 124.02 56.8 124.31 ;
      RECT  56.93 124.56 57.22 124.85 ;
      RECT  55.81 125.81 56.14 126.07 ;
      RECT  58.89 126.07 62.89 126.52 ;
      RECT  58.89 120.78 62.89 121.19 ;
      RECT  59.77 121.9 60.1 122.05 ;
      RECT  61.79 121.19 62.09 121.6 ;
      RECT  59.79 122.05 60.08 122.21 ;
      RECT  59.74 121.19 60.03 121.66 ;
      RECT  61.63 125.81 61.95 126.07 ;
      RECT  60.51 124.02 60.8 124.31 ;
      RECT  60.93 124.56 61.22 124.85 ;
      RECT  59.81 125.81 60.14 126.07 ;
      RECT  54.89 122.05 62.89 122.21 ;
      RECT  54.89 126.07 58.89 126.52 ;
      RECT  58.89 126.07 62.89 126.52 ;
      RECT  58.89 120.78 62.89 121.19 ;
      RECT  54.89 120.78 58.89 121.19 ;
      RECT  46.89 30.31 50.89 30.76 ;
      RECT  46.89 25.02 50.89 25.43 ;
      RECT  47.77 26.14 48.1 26.29 ;
      RECT  49.79 25.43 50.09 25.84 ;
      RECT  47.79 26.29 48.08 26.45 ;
      RECT  47.74 25.43 48.03 25.9 ;
      RECT  49.63 30.05 49.95 30.31 ;
      RECT  48.51 28.26 48.8 28.55 ;
      RECT  48.93 28.8 49.22 29.09 ;
      RECT  47.81 30.05 48.14 30.31 ;
      RECT  46.89 30.77 50.89 30.32 ;
      RECT  46.89 36.06 50.89 35.65 ;
      RECT  47.77 34.94 48.1 34.79 ;
      RECT  49.79 35.65 50.09 35.24 ;
      RECT  47.79 34.79 48.08 34.63 ;
      RECT  47.74 35.65 48.03 35.18 ;
      RECT  49.63 31.03 49.95 30.77 ;
      RECT  48.51 32.82 48.8 32.53 ;
      RECT  48.93 32.28 49.22 31.99 ;
      RECT  47.81 31.03 48.14 30.77 ;
      RECT  46.89 40.95 50.89 41.4 ;
      RECT  46.89 35.66 50.89 36.07 ;
      RECT  47.77 36.78 48.1 36.93 ;
      RECT  49.79 36.07 50.09 36.48 ;
      RECT  47.79 36.93 48.08 37.09 ;
      RECT  47.74 36.07 48.03 36.54 ;
      RECT  49.63 40.69 49.95 40.95 ;
      RECT  48.51 38.9 48.8 39.19 ;
      RECT  48.93 39.44 49.22 39.73 ;
      RECT  47.81 40.69 48.14 40.95 ;
      RECT  46.89 41.41 50.89 40.96 ;
      RECT  46.89 46.7 50.89 46.29 ;
      RECT  47.77 45.58 48.1 45.43 ;
      RECT  49.79 46.29 50.09 45.88 ;
      RECT  47.79 45.43 48.08 45.27 ;
      RECT  47.74 46.29 48.03 45.82 ;
      RECT  49.63 41.67 49.95 41.41 ;
      RECT  48.51 43.46 48.8 43.17 ;
      RECT  48.93 42.92 49.22 42.63 ;
      RECT  47.81 41.67 48.14 41.41 ;
      RECT  46.89 51.59 50.89 52.04 ;
      RECT  46.89 46.3 50.89 46.71 ;
      RECT  47.77 47.42 48.1 47.57 ;
      RECT  49.79 46.71 50.09 47.12 ;
      RECT  47.79 47.57 48.08 47.73 ;
      RECT  47.74 46.71 48.03 47.18 ;
      RECT  49.63 51.33 49.95 51.59 ;
      RECT  48.51 49.54 48.8 49.83 ;
      RECT  48.93 50.08 49.22 50.37 ;
      RECT  47.81 51.33 48.14 51.59 ;
      RECT  46.89 52.05 50.89 51.6 ;
      RECT  46.89 57.34 50.89 56.93 ;
      RECT  47.77 56.22 48.1 56.07 ;
      RECT  49.79 56.93 50.09 56.52 ;
      RECT  47.79 56.07 48.08 55.91 ;
      RECT  47.74 56.93 48.03 56.46 ;
      RECT  49.63 52.31 49.95 52.05 ;
      RECT  48.51 54.1 48.8 53.81 ;
      RECT  48.93 53.56 49.22 53.27 ;
      RECT  47.81 52.31 48.14 52.05 ;
      RECT  46.89 62.23 50.89 62.68 ;
      RECT  46.89 56.94 50.89 57.35 ;
      RECT  47.77 58.06 48.1 58.21 ;
      RECT  49.79 57.35 50.09 57.76 ;
      RECT  47.79 58.21 48.08 58.37 ;
      RECT  47.74 57.35 48.03 57.82 ;
      RECT  49.63 61.97 49.95 62.23 ;
      RECT  48.51 60.18 48.8 60.47 ;
      RECT  48.93 60.72 49.22 61.01 ;
      RECT  47.81 61.97 48.14 62.23 ;
      RECT  46.89 62.69 50.89 62.24 ;
      RECT  46.89 67.98 50.89 67.57 ;
      RECT  47.77 66.86 48.1 66.71 ;
      RECT  49.79 67.57 50.09 67.16 ;
      RECT  47.79 66.71 48.08 66.55 ;
      RECT  47.74 67.57 48.03 67.1 ;
      RECT  49.63 62.95 49.95 62.69 ;
      RECT  48.51 64.74 48.8 64.45 ;
      RECT  48.93 64.2 49.22 63.91 ;
      RECT  47.81 62.95 48.14 62.69 ;
      RECT  46.89 72.87 50.89 73.32 ;
      RECT  46.89 67.58 50.89 67.99 ;
      RECT  47.77 68.7 48.1 68.85 ;
      RECT  49.79 67.99 50.09 68.4 ;
      RECT  47.79 68.85 48.08 69.01 ;
      RECT  47.74 67.99 48.03 68.46 ;
      RECT  49.63 72.61 49.95 72.87 ;
      RECT  48.51 70.82 48.8 71.11 ;
      RECT  48.93 71.36 49.22 71.65 ;
      RECT  47.81 72.61 48.14 72.87 ;
      RECT  46.89 73.33 50.89 72.88 ;
      RECT  46.89 78.62 50.89 78.21 ;
      RECT  47.77 77.5 48.1 77.35 ;
      RECT  49.79 78.21 50.09 77.8 ;
      RECT  47.79 77.35 48.08 77.19 ;
      RECT  47.74 78.21 48.03 77.74 ;
      RECT  49.63 73.59 49.95 73.33 ;
      RECT  48.51 75.38 48.8 75.09 ;
      RECT  48.93 74.84 49.22 74.55 ;
      RECT  47.81 73.59 48.14 73.33 ;
      RECT  46.89 83.51 50.89 83.96 ;
      RECT  46.89 78.22 50.89 78.63 ;
      RECT  47.77 79.34 48.1 79.49 ;
      RECT  49.79 78.63 50.09 79.04 ;
      RECT  47.79 79.49 48.08 79.65 ;
      RECT  47.74 78.63 48.03 79.1 ;
      RECT  49.63 83.25 49.95 83.51 ;
      RECT  48.51 81.46 48.8 81.75 ;
      RECT  48.93 82.0 49.22 82.29 ;
      RECT  47.81 83.25 48.14 83.51 ;
      RECT  46.89 83.97 50.89 83.52 ;
      RECT  46.89 89.26 50.89 88.85 ;
      RECT  47.77 88.14 48.1 87.99 ;
      RECT  49.79 88.85 50.09 88.44 ;
      RECT  47.79 87.99 48.08 87.83 ;
      RECT  47.74 88.85 48.03 88.38 ;
      RECT  49.63 84.23 49.95 83.97 ;
      RECT  48.51 86.02 48.8 85.73 ;
      RECT  48.93 85.48 49.22 85.19 ;
      RECT  47.81 84.23 48.14 83.97 ;
      RECT  46.89 94.15 50.89 94.6 ;
      RECT  46.89 88.86 50.89 89.27 ;
      RECT  47.77 89.98 48.1 90.13 ;
      RECT  49.79 89.27 50.09 89.68 ;
      RECT  47.79 90.13 48.08 90.29 ;
      RECT  47.74 89.27 48.03 89.74 ;
      RECT  49.63 93.89 49.95 94.15 ;
      RECT  48.51 92.1 48.8 92.39 ;
      RECT  48.93 92.64 49.22 92.93 ;
      RECT  47.81 93.89 48.14 94.15 ;
      RECT  46.89 94.61 50.89 94.16 ;
      RECT  46.89 99.9 50.89 99.49 ;
      RECT  47.77 98.78 48.1 98.63 ;
      RECT  49.79 99.49 50.09 99.08 ;
      RECT  47.79 98.63 48.08 98.47 ;
      RECT  47.74 99.49 48.03 99.02 ;
      RECT  49.63 94.87 49.95 94.61 ;
      RECT  48.51 96.66 48.8 96.37 ;
      RECT  48.93 96.12 49.22 95.83 ;
      RECT  47.81 94.87 48.14 94.61 ;
      RECT  46.89 104.79 50.89 105.24 ;
      RECT  46.89 99.5 50.89 99.91 ;
      RECT  47.77 100.62 48.1 100.77 ;
      RECT  49.79 99.91 50.09 100.32 ;
      RECT  47.79 100.77 48.08 100.93 ;
      RECT  47.74 99.91 48.03 100.38 ;
      RECT  49.63 104.53 49.95 104.79 ;
      RECT  48.51 102.74 48.8 103.03 ;
      RECT  48.93 103.28 49.22 103.57 ;
      RECT  47.81 104.53 48.14 104.79 ;
      RECT  46.89 105.25 50.89 104.8 ;
      RECT  46.89 110.54 50.89 110.13 ;
      RECT  47.77 109.42 48.1 109.27 ;
      RECT  49.79 110.13 50.09 109.72 ;
      RECT  47.79 109.27 48.08 109.11 ;
      RECT  47.74 110.13 48.03 109.66 ;
      RECT  49.63 105.51 49.95 105.25 ;
      RECT  48.51 107.3 48.8 107.01 ;
      RECT  48.93 106.76 49.22 106.47 ;
      RECT  47.81 105.51 48.14 105.25 ;
      RECT  46.89 115.43 50.89 115.88 ;
      RECT  46.89 110.14 50.89 110.55 ;
      RECT  47.77 111.26 48.1 111.41 ;
      RECT  49.79 110.55 50.09 110.96 ;
      RECT  47.79 111.41 48.08 111.57 ;
      RECT  47.74 110.55 48.03 111.02 ;
      RECT  49.63 115.17 49.95 115.43 ;
      RECT  48.51 113.38 48.8 113.67 ;
      RECT  48.93 113.92 49.22 114.21 ;
      RECT  47.81 115.17 48.14 115.43 ;
      RECT  46.89 115.89 50.89 115.44 ;
      RECT  46.89 121.18 50.89 120.77 ;
      RECT  47.77 120.06 48.1 119.91 ;
      RECT  49.79 120.77 50.09 120.36 ;
      RECT  47.79 119.91 48.08 119.75 ;
      RECT  47.74 120.77 48.03 120.3 ;
      RECT  49.63 116.15 49.95 115.89 ;
      RECT  48.51 117.94 48.8 117.65 ;
      RECT  48.93 117.4 49.22 117.11 ;
      RECT  47.81 116.15 48.14 115.89 ;
      RECT  46.89 126.07 50.89 126.52 ;
      RECT  46.89 120.78 50.89 121.19 ;
      RECT  47.77 121.9 48.1 122.05 ;
      RECT  49.79 121.19 50.09 121.6 ;
      RECT  47.79 122.05 48.08 122.21 ;
      RECT  47.74 121.19 48.03 121.66 ;
      RECT  49.63 125.81 49.95 126.07 ;
      RECT  48.51 124.02 48.8 124.31 ;
      RECT  48.93 124.56 49.22 124.85 ;
      RECT  47.81 125.81 48.14 126.07 ;
      RECT  46.89 26.29 50.89 26.45 ;
      RECT  46.89 34.63 50.89 34.79 ;
      RECT  46.89 36.93 50.89 37.09 ;
      RECT  46.89 45.27 50.89 45.43 ;
      RECT  46.89 47.57 50.89 47.73 ;
      RECT  46.89 55.91 50.89 56.07 ;
      RECT  46.89 58.21 50.89 58.37 ;
      RECT  46.89 66.55 50.89 66.71 ;
      RECT  46.89 68.85 50.89 69.01 ;
      RECT  46.89 77.19 50.89 77.35 ;
      RECT  46.89 79.49 50.89 79.65 ;
      RECT  46.89 87.83 50.89 87.99 ;
      RECT  46.89 90.13 50.89 90.29 ;
      RECT  46.89 98.47 50.89 98.63 ;
      RECT  46.89 100.77 50.89 100.93 ;
      RECT  46.89 109.11 50.89 109.27 ;
      RECT  46.89 111.41 50.89 111.57 ;
      RECT  46.89 119.75 50.89 119.91 ;
      RECT  46.89 122.05 50.89 122.21 ;
      RECT  46.89 30.32 50.89 30.77 ;
      RECT  46.89 30.31 50.89 30.76 ;
      RECT  46.89 94.16 50.89 94.61 ;
      RECT  46.89 62.24 50.89 62.69 ;
      RECT  46.89 83.52 50.89 83.97 ;
      RECT  46.89 51.59 50.89 52.04 ;
      RECT  46.89 72.88 50.89 73.33 ;
      RECT  46.89 83.51 50.89 83.96 ;
      RECT  46.89 94.15 50.89 94.6 ;
      RECT  46.89 115.44 50.89 115.89 ;
      RECT  46.89 40.96 50.89 41.41 ;
      RECT  46.89 126.07 50.89 126.52 ;
      RECT  46.89 51.6 50.89 52.05 ;
      RECT  46.89 62.23 50.89 62.68 ;
      RECT  46.89 115.43 50.89 115.88 ;
      RECT  46.89 72.87 50.89 73.32 ;
      RECT  46.89 104.79 50.89 105.24 ;
      RECT  46.89 40.95 50.89 41.4 ;
      RECT  46.89 104.8 50.89 105.25 ;
      RECT  46.89 99.49 50.89 99.9 ;
      RECT  46.89 110.13 50.89 110.54 ;
      RECT  46.89 56.93 50.89 57.34 ;
      RECT  46.89 110.14 50.89 110.55 ;
      RECT  46.89 120.77 50.89 121.18 ;
      RECT  46.89 99.5 50.89 99.91 ;
      RECT  46.89 46.3 50.89 46.71 ;
      RECT  46.89 78.22 50.89 78.63 ;
      RECT  46.89 46.29 50.89 46.7 ;
      RECT  46.89 78.21 50.89 78.62 ;
      RECT  46.89 25.02 50.89 25.43 ;
      RECT  46.89 120.78 50.89 121.19 ;
      RECT  46.89 88.86 50.89 89.27 ;
      RECT  46.89 67.58 50.89 67.99 ;
      RECT  46.89 56.94 50.89 57.35 ;
      RECT  46.89 67.57 50.89 67.98 ;
      RECT  46.89 35.66 50.89 36.07 ;
      RECT  46.89 88.85 50.89 89.26 ;
      RECT  46.89 35.65 50.89 36.06 ;
      RECT  62.89 30.31 66.89 30.76 ;
      RECT  62.89 25.02 66.89 25.43 ;
      RECT  63.77 26.14 64.1 26.29 ;
      RECT  65.79 25.43 66.09 25.84 ;
      RECT  63.79 26.29 64.08 26.45 ;
      RECT  63.74 25.43 64.03 25.9 ;
      RECT  65.63 30.05 65.95 30.31 ;
      RECT  64.51 28.26 64.8 28.55 ;
      RECT  64.93 28.8 65.22 29.09 ;
      RECT  63.81 30.05 64.14 30.31 ;
      RECT  62.89 30.77 66.89 30.32 ;
      RECT  62.89 36.06 66.89 35.65 ;
      RECT  63.77 34.94 64.1 34.79 ;
      RECT  65.79 35.65 66.09 35.24 ;
      RECT  63.79 34.79 64.08 34.63 ;
      RECT  63.74 35.65 64.03 35.18 ;
      RECT  65.63 31.03 65.95 30.77 ;
      RECT  64.51 32.82 64.8 32.53 ;
      RECT  64.93 32.28 65.22 31.99 ;
      RECT  63.81 31.03 64.14 30.77 ;
      RECT  62.89 40.95 66.89 41.4 ;
      RECT  62.89 35.66 66.89 36.07 ;
      RECT  63.77 36.78 64.1 36.93 ;
      RECT  65.79 36.07 66.09 36.48 ;
      RECT  63.79 36.93 64.08 37.09 ;
      RECT  63.74 36.07 64.03 36.54 ;
      RECT  65.63 40.69 65.95 40.95 ;
      RECT  64.51 38.9 64.8 39.19 ;
      RECT  64.93 39.44 65.22 39.73 ;
      RECT  63.81 40.69 64.14 40.95 ;
      RECT  62.89 41.41 66.89 40.96 ;
      RECT  62.89 46.7 66.89 46.29 ;
      RECT  63.77 45.58 64.1 45.43 ;
      RECT  65.79 46.29 66.09 45.88 ;
      RECT  63.79 45.43 64.08 45.27 ;
      RECT  63.74 46.29 64.03 45.82 ;
      RECT  65.63 41.67 65.95 41.41 ;
      RECT  64.51 43.46 64.8 43.17 ;
      RECT  64.93 42.92 65.22 42.63 ;
      RECT  63.81 41.67 64.14 41.41 ;
      RECT  62.89 51.59 66.89 52.04 ;
      RECT  62.89 46.3 66.89 46.71 ;
      RECT  63.77 47.42 64.1 47.57 ;
      RECT  65.79 46.71 66.09 47.12 ;
      RECT  63.79 47.57 64.08 47.73 ;
      RECT  63.74 46.71 64.03 47.18 ;
      RECT  65.63 51.33 65.95 51.59 ;
      RECT  64.51 49.54 64.8 49.83 ;
      RECT  64.93 50.08 65.22 50.37 ;
      RECT  63.81 51.33 64.14 51.59 ;
      RECT  62.89 52.05 66.89 51.6 ;
      RECT  62.89 57.34 66.89 56.93 ;
      RECT  63.77 56.22 64.1 56.07 ;
      RECT  65.79 56.93 66.09 56.52 ;
      RECT  63.79 56.07 64.08 55.91 ;
      RECT  63.74 56.93 64.03 56.46 ;
      RECT  65.63 52.31 65.95 52.05 ;
      RECT  64.51 54.1 64.8 53.81 ;
      RECT  64.93 53.56 65.22 53.27 ;
      RECT  63.81 52.31 64.14 52.05 ;
      RECT  62.89 62.23 66.89 62.68 ;
      RECT  62.89 56.94 66.89 57.35 ;
      RECT  63.77 58.06 64.1 58.21 ;
      RECT  65.79 57.35 66.09 57.76 ;
      RECT  63.79 58.21 64.08 58.37 ;
      RECT  63.74 57.35 64.03 57.82 ;
      RECT  65.63 61.97 65.95 62.23 ;
      RECT  64.51 60.18 64.8 60.47 ;
      RECT  64.93 60.72 65.22 61.01 ;
      RECT  63.81 61.97 64.14 62.23 ;
      RECT  62.89 62.69 66.89 62.24 ;
      RECT  62.89 67.98 66.89 67.57 ;
      RECT  63.77 66.86 64.1 66.71 ;
      RECT  65.79 67.57 66.09 67.16 ;
      RECT  63.79 66.71 64.08 66.55 ;
      RECT  63.74 67.57 64.03 67.1 ;
      RECT  65.63 62.95 65.95 62.69 ;
      RECT  64.51 64.74 64.8 64.45 ;
      RECT  64.93 64.2 65.22 63.91 ;
      RECT  63.81 62.95 64.14 62.69 ;
      RECT  62.89 72.87 66.89 73.32 ;
      RECT  62.89 67.58 66.89 67.99 ;
      RECT  63.77 68.7 64.1 68.85 ;
      RECT  65.79 67.99 66.09 68.4 ;
      RECT  63.79 68.85 64.08 69.01 ;
      RECT  63.74 67.99 64.03 68.46 ;
      RECT  65.63 72.61 65.95 72.87 ;
      RECT  64.51 70.82 64.8 71.11 ;
      RECT  64.93 71.36 65.22 71.65 ;
      RECT  63.81 72.61 64.14 72.87 ;
      RECT  62.89 73.33 66.89 72.88 ;
      RECT  62.89 78.62 66.89 78.21 ;
      RECT  63.77 77.5 64.1 77.35 ;
      RECT  65.79 78.21 66.09 77.8 ;
      RECT  63.79 77.35 64.08 77.19 ;
      RECT  63.74 78.21 64.03 77.74 ;
      RECT  65.63 73.59 65.95 73.33 ;
      RECT  64.51 75.38 64.8 75.09 ;
      RECT  64.93 74.84 65.22 74.55 ;
      RECT  63.81 73.59 64.14 73.33 ;
      RECT  62.89 83.51 66.89 83.96 ;
      RECT  62.89 78.22 66.89 78.63 ;
      RECT  63.77 79.34 64.1 79.49 ;
      RECT  65.79 78.63 66.09 79.04 ;
      RECT  63.79 79.49 64.08 79.65 ;
      RECT  63.74 78.63 64.03 79.1 ;
      RECT  65.63 83.25 65.95 83.51 ;
      RECT  64.51 81.46 64.8 81.75 ;
      RECT  64.93 82.0 65.22 82.29 ;
      RECT  63.81 83.25 64.14 83.51 ;
      RECT  62.89 83.97 66.89 83.52 ;
      RECT  62.89 89.26 66.89 88.85 ;
      RECT  63.77 88.14 64.1 87.99 ;
      RECT  65.79 88.85 66.09 88.44 ;
      RECT  63.79 87.99 64.08 87.83 ;
      RECT  63.74 88.85 64.03 88.38 ;
      RECT  65.63 84.23 65.95 83.97 ;
      RECT  64.51 86.02 64.8 85.73 ;
      RECT  64.93 85.48 65.22 85.19 ;
      RECT  63.81 84.23 64.14 83.97 ;
      RECT  62.89 94.15 66.89 94.6 ;
      RECT  62.89 88.86 66.89 89.27 ;
      RECT  63.77 89.98 64.1 90.13 ;
      RECT  65.79 89.27 66.09 89.68 ;
      RECT  63.79 90.13 64.08 90.29 ;
      RECT  63.74 89.27 64.03 89.74 ;
      RECT  65.63 93.89 65.95 94.15 ;
      RECT  64.51 92.1 64.8 92.39 ;
      RECT  64.93 92.64 65.22 92.93 ;
      RECT  63.81 93.89 64.14 94.15 ;
      RECT  62.89 94.61 66.89 94.16 ;
      RECT  62.89 99.9 66.89 99.49 ;
      RECT  63.77 98.78 64.1 98.63 ;
      RECT  65.79 99.49 66.09 99.08 ;
      RECT  63.79 98.63 64.08 98.47 ;
      RECT  63.74 99.49 64.03 99.02 ;
      RECT  65.63 94.87 65.95 94.61 ;
      RECT  64.51 96.66 64.8 96.37 ;
      RECT  64.93 96.12 65.22 95.83 ;
      RECT  63.81 94.87 64.14 94.61 ;
      RECT  62.89 104.79 66.89 105.24 ;
      RECT  62.89 99.5 66.89 99.91 ;
      RECT  63.77 100.62 64.1 100.77 ;
      RECT  65.79 99.91 66.09 100.32 ;
      RECT  63.79 100.77 64.08 100.93 ;
      RECT  63.74 99.91 64.03 100.38 ;
      RECT  65.63 104.53 65.95 104.79 ;
      RECT  64.51 102.74 64.8 103.03 ;
      RECT  64.93 103.28 65.22 103.57 ;
      RECT  63.81 104.53 64.14 104.79 ;
      RECT  62.89 105.25 66.89 104.8 ;
      RECT  62.89 110.54 66.89 110.13 ;
      RECT  63.77 109.42 64.1 109.27 ;
      RECT  65.79 110.13 66.09 109.72 ;
      RECT  63.79 109.27 64.08 109.11 ;
      RECT  63.74 110.13 64.03 109.66 ;
      RECT  65.63 105.51 65.95 105.25 ;
      RECT  64.51 107.3 64.8 107.01 ;
      RECT  64.93 106.76 65.22 106.47 ;
      RECT  63.81 105.51 64.14 105.25 ;
      RECT  62.89 115.43 66.89 115.88 ;
      RECT  62.89 110.14 66.89 110.55 ;
      RECT  63.77 111.26 64.1 111.41 ;
      RECT  65.79 110.55 66.09 110.96 ;
      RECT  63.79 111.41 64.08 111.57 ;
      RECT  63.74 110.55 64.03 111.02 ;
      RECT  65.63 115.17 65.95 115.43 ;
      RECT  64.51 113.38 64.8 113.67 ;
      RECT  64.93 113.92 65.22 114.21 ;
      RECT  63.81 115.17 64.14 115.43 ;
      RECT  62.89 115.89 66.89 115.44 ;
      RECT  62.89 121.18 66.89 120.77 ;
      RECT  63.77 120.06 64.1 119.91 ;
      RECT  65.79 120.77 66.09 120.36 ;
      RECT  63.79 119.91 64.08 119.75 ;
      RECT  63.74 120.77 64.03 120.3 ;
      RECT  65.63 116.15 65.95 115.89 ;
      RECT  64.51 117.94 64.8 117.65 ;
      RECT  64.93 117.4 65.22 117.11 ;
      RECT  63.81 116.15 64.14 115.89 ;
      RECT  62.89 126.07 66.89 126.52 ;
      RECT  62.89 120.78 66.89 121.19 ;
      RECT  63.77 121.9 64.1 122.05 ;
      RECT  65.79 121.19 66.09 121.6 ;
      RECT  63.79 122.05 64.08 122.21 ;
      RECT  63.74 121.19 64.03 121.66 ;
      RECT  65.63 125.81 65.95 126.07 ;
      RECT  64.51 124.02 64.8 124.31 ;
      RECT  64.93 124.56 65.22 124.85 ;
      RECT  63.81 125.81 64.14 126.07 ;
      RECT  62.89 26.29 66.89 26.45 ;
      RECT  62.89 34.63 66.89 34.79 ;
      RECT  62.89 36.93 66.89 37.09 ;
      RECT  62.89 45.27 66.89 45.43 ;
      RECT  62.89 47.57 66.89 47.73 ;
      RECT  62.89 55.91 66.89 56.07 ;
      RECT  62.89 58.21 66.89 58.37 ;
      RECT  62.89 66.55 66.89 66.71 ;
      RECT  62.89 68.85 66.89 69.01 ;
      RECT  62.89 77.19 66.89 77.35 ;
      RECT  62.89 79.49 66.89 79.65 ;
      RECT  62.89 87.83 66.89 87.99 ;
      RECT  62.89 90.13 66.89 90.29 ;
      RECT  62.89 98.47 66.89 98.63 ;
      RECT  62.89 100.77 66.89 100.93 ;
      RECT  62.89 109.11 66.89 109.27 ;
      RECT  62.89 111.41 66.89 111.57 ;
      RECT  62.89 119.75 66.89 119.91 ;
      RECT  62.89 122.05 66.89 122.21 ;
      RECT  62.89 30.32 66.89 30.77 ;
      RECT  62.89 30.31 66.89 30.76 ;
      RECT  62.89 94.16 66.89 94.61 ;
      RECT  62.89 62.24 66.89 62.69 ;
      RECT  62.89 83.52 66.89 83.97 ;
      RECT  62.89 51.59 66.89 52.04 ;
      RECT  62.89 72.88 66.89 73.33 ;
      RECT  62.89 83.51 66.89 83.96 ;
      RECT  62.89 94.15 66.89 94.6 ;
      RECT  62.89 115.44 66.89 115.89 ;
      RECT  62.89 40.96 66.89 41.41 ;
      RECT  62.89 126.07 66.89 126.52 ;
      RECT  62.89 51.6 66.89 52.05 ;
      RECT  62.89 62.23 66.89 62.68 ;
      RECT  62.89 115.43 66.89 115.88 ;
      RECT  62.89 72.87 66.89 73.32 ;
      RECT  62.89 104.79 66.89 105.24 ;
      RECT  62.89 40.95 66.89 41.4 ;
      RECT  62.89 104.8 66.89 105.25 ;
      RECT  62.89 99.49 66.89 99.9 ;
      RECT  62.89 110.13 66.89 110.54 ;
      RECT  62.89 56.93 66.89 57.34 ;
      RECT  62.89 110.14 66.89 110.55 ;
      RECT  62.89 120.77 66.89 121.18 ;
      RECT  62.89 99.5 66.89 99.91 ;
      RECT  62.89 46.3 66.89 46.71 ;
      RECT  62.89 78.22 66.89 78.63 ;
      RECT  62.89 46.29 66.89 46.7 ;
      RECT  62.89 78.21 66.89 78.62 ;
      RECT  62.89 25.02 66.89 25.43 ;
      RECT  62.89 120.78 66.89 121.19 ;
      RECT  62.89 88.86 66.89 89.27 ;
      RECT  62.89 67.58 66.89 67.99 ;
      RECT  62.89 56.94 66.89 57.35 ;
      RECT  62.89 67.57 66.89 67.98 ;
      RECT  62.89 35.66 66.89 36.07 ;
      RECT  62.89 88.85 66.89 89.26 ;
      RECT  62.89 35.65 66.89 36.06 ;
      RECT  45.99 34.63 67.79 34.79 ;
      RECT  45.99 36.93 67.79 37.09 ;
      RECT  45.99 45.27 67.79 45.43 ;
      RECT  45.99 47.57 67.79 47.73 ;
      RECT  45.99 55.91 67.79 56.07 ;
      RECT  45.99 58.21 67.79 58.37 ;
      RECT  45.99 66.55 67.79 66.71 ;
      RECT  45.99 68.85 67.79 69.01 ;
      RECT  45.99 77.19 67.79 77.35 ;
      RECT  45.99 79.49 67.79 79.65 ;
      RECT  45.99 87.83 67.79 87.99 ;
      RECT  45.99 90.13 67.79 90.29 ;
      RECT  45.99 98.47 67.79 98.63 ;
      RECT  45.99 100.77 67.79 100.93 ;
      RECT  45.99 109.11 67.79 109.27 ;
      RECT  45.99 111.41 67.79 111.57 ;
      RECT  45.99 119.75 67.79 119.91 ;
      RECT  50.89 62.24 54.89 62.69 ;
      RECT  50.89 51.59 54.89 52.04 ;
      RECT  50.89 83.52 54.89 83.97 ;
      RECT  50.89 40.95 54.89 41.4 ;
      RECT  50.89 51.6 54.89 52.05 ;
      RECT  50.89 40.96 54.89 41.41 ;
      RECT  50.89 62.23 54.89 62.68 ;
      RECT  50.89 115.44 54.89 115.89 ;
      RECT  50.89 72.88 54.89 73.33 ;
      RECT  50.89 94.16 54.89 94.61 ;
      RECT  50.89 115.43 54.89 115.88 ;
      RECT  50.89 104.79 54.89 105.24 ;
      RECT  50.89 104.8 54.89 105.25 ;
      RECT  50.89 83.51 54.89 83.96 ;
      RECT  50.89 72.87 54.89 73.32 ;
      RECT  50.89 30.32 54.89 30.77 ;
      RECT  50.89 94.15 54.89 94.6 ;
      RECT  50.89 110.13 54.89 110.54 ;
      RECT  50.89 35.65 54.89 36.06 ;
      RECT  50.89 120.77 54.89 121.18 ;
      RECT  50.89 78.22 54.89 78.63 ;
      RECT  50.89 56.94 54.89 57.35 ;
      RECT  50.89 78.21 54.89 78.62 ;
      RECT  50.89 88.85 54.89 89.26 ;
      RECT  50.89 46.29 54.89 46.7 ;
      RECT  50.89 88.86 54.89 89.27 ;
      RECT  50.89 67.58 54.89 67.99 ;
      RECT  50.89 67.57 54.89 67.98 ;
      RECT  50.89 99.49 54.89 99.9 ;
      RECT  50.89 110.14 54.89 110.55 ;
      RECT  50.89 56.93 54.89 57.34 ;
      RECT  50.89 99.5 54.89 99.91 ;
      RECT  50.89 46.3 54.89 46.71 ;
      RECT  50.89 35.66 54.89 36.07 ;
      RECT  50.89 17.14 54.89 17.28 ;
      RECT  54.89 17.14 58.89 17.28 ;
      RECT  58.89 17.14 62.89 17.28 ;
      RECT  45.99 17.14 62.89 17.28 ;
      RECT  54.89 10.26 58.89 10.4 ;
      RECT  56.32 10.02 56.61 10.11 ;
      RECT  57.63 10.61 57.96 10.94 ;
      RECT  56.39 11.23 56.72 11.56 ;
      RECT  55.25 12.39 55.54 12.48 ;
      RECT  55.15 11.06 55.44 11.11 ;
      RECT  55.15 10.82 55.46 11.06 ;
      RECT  54.89 12.25 58.89 12.39 ;
      RECT  57.49 9.82 57.78 9.88 ;
      RECT  56.32 9.88 57.78 10.02 ;
      RECT  55.25 12.19 55.54 12.25 ;
      RECT  57.49 10.02 57.78 10.11 ;
      RECT  55.32 10.4 55.46 10.82 ;
      RECT  54.89 9.12 58.89 9.41 ;
      RECT  54.89 13.58 58.89 13.87 ;
      RECT  56.32 9.82 56.61 9.88 ;
      RECT  58.89 10.26 62.89 10.4 ;
      RECT  60.32 10.02 60.61 10.11 ;
      RECT  61.63 10.61 61.96 10.94 ;
      RECT  60.39 11.23 60.72 11.56 ;
      RECT  59.25 12.39 59.54 12.48 ;
      RECT  59.15 11.06 59.44 11.11 ;
      RECT  59.15 10.82 59.46 11.06 ;
      RECT  58.89 12.25 62.89 12.39 ;
      RECT  61.49 9.82 61.78 9.88 ;
      RECT  60.32 9.88 61.78 10.02 ;
      RECT  59.25 12.19 59.54 12.25 ;
      RECT  61.49 10.02 61.78 10.11 ;
      RECT  59.32 10.4 59.46 10.82 ;
      RECT  58.89 9.12 62.89 9.41 ;
      RECT  58.89 13.58 62.89 13.87 ;
      RECT  60.32 9.82 60.61 9.88 ;
      RECT  54.89 12.25 58.89 12.39 ;
      RECT  58.89 12.25 62.89 12.39 ;
      RECT  45.99 10.87 62.89 11.01 ;
      RECT  57.66 3.55 57.96 3.6 ;
      RECT  56.06 6.94 68.3 7.39 ;
      RECT  57.66 3.8 57.96 3.85 ;
      RECT  65.83 3.97 66.16 4.01 ;
      RECT  59.97 3.08 60.27 5.7 ;
      RECT  66.28 5.41 66.58 5.7 ;
      RECT  56.06 1.15 68.3 1.57 ;
      RECT  66.32 3.37 66.58 5.41 ;
      RECT  66.28 3.08 66.58 3.37 ;
      RECT  67.83 4.41 68.13 4.7 ;
      RECT  67.99 3.04 68.29 3.33 ;
      RECT  56.06 3.6 57.96 3.8 ;
      RECT  56.16 3.02 56.49 3.35 ;
      RECT  61.22 3.68 66.16 3.97 ;
      RECT  61.67 4.41 65.5 4.7 ;
      RECT  61.66 3.55 61.96 3.6 ;
      RECT  60.06 6.94 72.3 7.39 ;
      RECT  61.66 3.8 61.96 3.85 ;
      RECT  69.83 3.97 70.16 4.01 ;
      RECT  63.97 3.08 64.27 5.7 ;
      RECT  70.28 5.41 70.58 5.7 ;
      RECT  60.06 1.15 72.3 1.57 ;
      RECT  70.32 3.37 70.58 5.41 ;
      RECT  70.28 3.08 70.58 3.37 ;
      RECT  71.83 4.41 72.13 4.7 ;
      RECT  71.99 3.04 72.29 3.33 ;
      RECT  60.06 3.6 61.96 3.8 ;
      RECT  60.16 3.02 60.49 3.35 ;
      RECT  65.22 3.68 70.16 3.97 ;
      RECT  65.67 4.41 69.5 4.7 ;
      RECT  45.99 3.68 72.3 3.82 ;
      RECT  54.89 12.39 58.89 12.25 ;
      RECT  58.89 12.39 62.89 12.25 ;
      RECT  45.99 11.01 62.89 10.87 ;
      RECT  45.99 17.28 62.89 17.14 ;
      RECT  45.99 3.82 72.3 3.68 ;
      RECT  54.89 12.25 58.89 12.39 ;
      RECT  58.89 12.25 62.89 12.39 ;
      RECT  -45.26 -6.25 -44.73 -6.02 ;
      RECT  -49.48 -7.41 -49.15 -7.29 ;
      RECT  -44.76 -8.27 -44.56 -8.11 ;
      RECT  -46.91 -8.31 -46.58 -8.29 ;
      RECT  -52.59 -8.52 -52.28 -8.2 ;
      RECT  -52.84 -6.02 -39.71 -5.57 ;
      RECT  -50.6 -8.31 -50.27 -8.23 ;
      RECT  -49.48 -7.62 -49.15 -7.61 ;
      RECT  -50.56 -8.23 -50.36 -7.61 ;
      RECT  -48.02 -6.25 -47.49 -6.02 ;
      RECT  -45.4 -7.62 -45.07 -7.61 ;
      RECT  -51.1 -7.28 -50.76 -6.96 ;
      RECT  -45.4 -7.41 -45.07 -7.29 ;
      RECT  -40.62 -6.25 -40.09 -6.02 ;
      RECT  -52.84 -10.26 -39.71 -9.85 ;
      RECT  -51.72 -8.51 -50.27 -8.31 ;
      RECT  -50.56 -7.61 -45.07 -7.41 ;
      RECT  -51.21 -9.85 -50.8 -9.48 ;
      RECT  -49.06 -9.85 -48.65 -9.48 ;
      RECT  -49.48 -8.11 -44.56 -7.86 ;
      RECT  -50.01 -8.31 -49.71 -8.25 ;
      RECT  -41.97 -6.25 -41.44 -6.02 ;
      RECT  -43.74 -6.25 -43.21 -6.02 ;
      RECT  -43.26 -9.85 -42.85 -9.48 ;
      RECT  -43.68 -7.62 -43.35 -7.61 ;
      RECT  -43.68 -7.41 -43.35 -7.29 ;
      RECT  -44.21 -8.51 -40.54 -8.31 ;
      RECT  -51.72 -8.31 -51.43 -8.25 ;
      RECT  -50.17 -9.85 -49.76 -9.48 ;
      RECT  -44.21 -8.31 -43.91 -8.27 ;
      RECT  -44.76 -7.61 -43.35 -7.41 ;
      RECT  -46.91 -8.62 -46.58 -8.52 ;
      RECT  -49.48 -7.86 -49.15 -7.83 ;
      RECT  -40.88 -8.61 -40.54 -8.51 ;
      RECT  -44.37 -9.85 -43.96 -9.48 ;
      RECT  -42.54 -7.96 -41.91 -7.64 ;
      RECT  -49.54 -6.25 -49.01 -6.02 ;
      RECT  -44.8 -8.6 -44.47 -8.27 ;
      RECT  -49.48 -8.16 -49.15 -8.11 ;
      RECT  -42.16 -9.85 -41.75 -9.48 ;
      RECT  -50.01 -8.52 -46.58 -8.31 ;
      RECT  -50.01 -8.56 -49.71 -8.52 ;
      RECT  -40.88 -8.31 -40.54 -8.28 ;
      RECT  -51.06 -6.25 -50.53 -6.02 ;
      RECT  -50.6 -8.56 -50.27 -8.51 ;
      RECT  -45.41 -9.85 -45.0 -9.48 ;
      RECT  -44.76 -7.86 -44.56 -7.61 ;
      RECT  -51.72 -8.54 -51.43 -8.51 ;
      RECT  -44.21 -8.58 -43.91 -8.51 ;
      RECT  -52.84 -6.02 -28.69 -5.57 ;
      RECT  -52.84 -10.26 -28.69 -9.81 ;
      RECT  -45.26 -5.35 -44.73 -5.58 ;
      RECT  -49.48 -4.19 -49.15 -4.31 ;
      RECT  -44.76 -3.33 -44.56 -3.49 ;
      RECT  -46.91 -3.29 -46.58 -3.31 ;
      RECT  -52.59 -3.08 -52.28 -3.4 ;
      RECT  -52.84 -5.58 -39.71 -6.03 ;
      RECT  -50.6 -3.29 -50.27 -3.37 ;
      RECT  -49.48 -3.98 -49.15 -3.99 ;
      RECT  -50.56 -3.37 -50.36 -3.99 ;
      RECT  -48.02 -5.35 -47.49 -5.58 ;
      RECT  -45.4 -3.98 -45.07 -3.99 ;
      RECT  -51.1 -4.32 -50.76 -4.64 ;
      RECT  -45.4 -4.19 -45.07 -4.31 ;
      RECT  -40.62 -5.35 -40.09 -5.58 ;
      RECT  -52.84 -1.34 -39.71 -1.75 ;
      RECT  -51.72 -3.09 -50.27 -3.29 ;
      RECT  -50.56 -3.99 -45.07 -4.19 ;
      RECT  -51.21 -1.75 -50.8 -2.12 ;
      RECT  -49.06 -1.75 -48.65 -2.12 ;
      RECT  -49.48 -3.49 -44.56 -3.74 ;
      RECT  -50.01 -3.29 -49.71 -3.35 ;
      RECT  -41.97 -5.35 -41.44 -5.58 ;
      RECT  -43.74 -5.35 -43.21 -5.58 ;
      RECT  -43.26 -1.75 -42.85 -2.12 ;
      RECT  -43.68 -3.98 -43.35 -3.99 ;
      RECT  -43.68 -4.19 -43.35 -4.31 ;
      RECT  -44.21 -3.09 -40.54 -3.29 ;
      RECT  -51.72 -3.29 -51.43 -3.35 ;
      RECT  -50.17 -1.75 -49.76 -2.12 ;
      RECT  -44.21 -3.29 -43.91 -3.33 ;
      RECT  -44.76 -3.99 -43.35 -4.19 ;
      RECT  -46.91 -2.98 -46.58 -3.08 ;
      RECT  -49.48 -3.74 -49.15 -3.77 ;
      RECT  -40.88 -2.99 -40.54 -3.09 ;
      RECT  -44.37 -1.75 -43.96 -2.12 ;
      RECT  -42.54 -3.64 -41.91 -3.96 ;
      RECT  -49.54 -5.35 -49.01 -5.58 ;
      RECT  -44.8 -3.0 -44.47 -3.33 ;
      RECT  -49.48 -3.44 -49.15 -3.49 ;
      RECT  -42.16 -1.75 -41.75 -2.12 ;
      RECT  -50.01 -3.08 -46.58 -3.29 ;
      RECT  -50.01 -3.04 -49.71 -3.08 ;
      RECT  -40.88 -3.29 -40.54 -3.32 ;
      RECT  -51.06 -5.35 -50.53 -5.58 ;
      RECT  -50.6 -3.04 -50.27 -3.09 ;
      RECT  -45.41 -1.75 -45.0 -2.12 ;
      RECT  -44.76 -3.74 -44.56 -3.99 ;
      RECT  -51.72 -3.06 -51.43 -3.09 ;
      RECT  -44.21 -3.02 -43.91 -3.09 ;
      RECT  -52.84 -5.58 -28.69 -6.03 ;
      RECT  -52.84 -1.34 -28.69 -1.79 ;
      RECT  -6.95 105.83 -6.42 106.06 ;
      RECT  -11.17 104.67 -10.84 104.79 ;
      RECT  -6.45 103.81 -6.25 103.97 ;
      RECT  -8.6 103.77 -8.27 103.79 ;
      RECT  -14.28 103.56 -13.97 103.88 ;
      RECT  -14.53 106.06 -1.4 106.51 ;
      RECT  -12.29 103.77 -11.96 103.85 ;
      RECT  -11.17 104.46 -10.84 104.47 ;
      RECT  -12.25 103.85 -12.05 104.47 ;
      RECT  -9.71 105.83 -9.18 106.06 ;
      RECT  -7.09 104.46 -6.76 104.47 ;
      RECT  -12.79 104.8 -12.45 105.12 ;
      RECT  -7.09 104.67 -6.76 104.79 ;
      RECT  -2.31 105.83 -1.78 106.06 ;
      RECT  -14.53 101.82 -1.4 102.23 ;
      RECT  -13.41 103.57 -11.96 103.77 ;
      RECT  -12.25 104.47 -6.76 104.67 ;
      RECT  -12.9 102.23 -12.49 102.6 ;
      RECT  -10.75 102.23 -10.34 102.6 ;
      RECT  -11.17 103.97 -6.25 104.22 ;
      RECT  -11.7 103.77 -11.4 103.83 ;
      RECT  -3.66 105.83 -3.13 106.06 ;
      RECT  -5.43 105.83 -4.9 106.06 ;
      RECT  -4.95 102.23 -4.54 102.6 ;
      RECT  -5.37 104.46 -5.04 104.47 ;
      RECT  -5.37 104.67 -5.04 104.79 ;
      RECT  -5.9 103.57 -2.23 103.77 ;
      RECT  -13.41 103.77 -13.12 103.83 ;
      RECT  -11.86 102.23 -11.45 102.6 ;
      RECT  -5.9 103.77 -5.6 103.81 ;
      RECT  -6.45 104.47 -5.04 104.67 ;
      RECT  -8.6 103.46 -8.27 103.56 ;
      RECT  -11.17 104.22 -10.84 104.25 ;
      RECT  -2.57 103.47 -2.23 103.57 ;
      RECT  -6.06 102.23 -5.65 102.6 ;
      RECT  -4.23 104.12 -3.6 104.44 ;
      RECT  -11.23 105.83 -10.7 106.06 ;
      RECT  -6.49 103.48 -6.16 103.81 ;
      RECT  -11.17 103.92 -10.84 103.97 ;
      RECT  -3.85 102.23 -3.44 102.6 ;
      RECT  -11.7 103.56 -8.27 103.77 ;
      RECT  -11.7 103.52 -11.4 103.56 ;
      RECT  -2.57 103.77 -2.23 103.8 ;
      RECT  -12.75 105.83 -12.22 106.06 ;
      RECT  -12.29 103.52 -11.96 103.57 ;
      RECT  -7.1 102.23 -6.69 102.6 ;
      RECT  -6.45 104.22 -6.25 104.47 ;
      RECT  -13.41 103.54 -13.12 103.57 ;
      RECT  -5.9 103.5 -5.6 103.57 ;
      RECT  -6.95 106.73 -6.42 106.5 ;
      RECT  -11.17 107.89 -10.84 107.77 ;
      RECT  -6.45 108.75 -6.25 108.59 ;
      RECT  -8.6 108.79 -8.27 108.77 ;
      RECT  -14.28 109.0 -13.97 108.68 ;
      RECT  -14.53 106.5 -1.4 106.05 ;
      RECT  -12.29 108.79 -11.96 108.71 ;
      RECT  -11.17 108.1 -10.84 108.09 ;
      RECT  -12.25 108.71 -12.05 108.09 ;
      RECT  -9.71 106.73 -9.18 106.5 ;
      RECT  -7.09 108.1 -6.76 108.09 ;
      RECT  -12.79 107.76 -12.45 107.44 ;
      RECT  -7.09 107.89 -6.76 107.77 ;
      RECT  -2.31 106.73 -1.78 106.5 ;
      RECT  -14.53 110.74 -1.4 110.33 ;
      RECT  -13.41 108.99 -11.96 108.79 ;
      RECT  -12.25 108.09 -6.76 107.89 ;
      RECT  -12.9 110.33 -12.49 109.96 ;
      RECT  -10.75 110.33 -10.34 109.96 ;
      RECT  -11.17 108.59 -6.25 108.34 ;
      RECT  -11.7 108.79 -11.4 108.73 ;
      RECT  -3.66 106.73 -3.13 106.5 ;
      RECT  -5.43 106.73 -4.9 106.5 ;
      RECT  -4.95 110.33 -4.54 109.96 ;
      RECT  -5.37 108.1 -5.04 108.09 ;
      RECT  -5.37 107.89 -5.04 107.77 ;
      RECT  -5.9 108.99 -2.23 108.79 ;
      RECT  -13.41 108.79 -13.12 108.73 ;
      RECT  -11.86 110.33 -11.45 109.96 ;
      RECT  -5.9 108.79 -5.6 108.75 ;
      RECT  -6.45 108.09 -5.04 107.89 ;
      RECT  -8.6 109.1 -8.27 109.0 ;
      RECT  -11.17 108.34 -10.84 108.31 ;
      RECT  -2.57 109.09 -2.23 108.99 ;
      RECT  -6.06 110.33 -5.65 109.96 ;
      RECT  -4.23 108.44 -3.6 108.12 ;
      RECT  -11.23 106.73 -10.7 106.5 ;
      RECT  -6.49 109.08 -6.16 108.75 ;
      RECT  -11.17 108.64 -10.84 108.59 ;
      RECT  -3.85 110.33 -3.44 109.96 ;
      RECT  -11.7 109.0 -8.27 108.79 ;
      RECT  -11.7 109.04 -11.4 109.0 ;
      RECT  -2.57 108.79 -2.23 108.76 ;
      RECT  -12.75 106.73 -12.22 106.5 ;
      RECT  -12.29 109.04 -11.96 108.99 ;
      RECT  -7.1 110.33 -6.69 109.96 ;
      RECT  -6.45 108.34 -6.25 108.09 ;
      RECT  -13.41 109.02 -13.12 108.99 ;
      RECT  -5.9 109.06 -5.6 108.99 ;
      RECT  -6.95 114.35 -6.42 114.58 ;
      RECT  -11.17 113.19 -10.84 113.31 ;
      RECT  -6.45 112.33 -6.25 112.49 ;
      RECT  -8.6 112.29 -8.27 112.31 ;
      RECT  -14.28 112.08 -13.97 112.4 ;
      RECT  -14.53 114.58 -1.4 115.03 ;
      RECT  -12.29 112.29 -11.96 112.37 ;
      RECT  -11.17 112.98 -10.84 112.99 ;
      RECT  -12.25 112.37 -12.05 112.99 ;
      RECT  -9.71 114.35 -9.18 114.58 ;
      RECT  -7.09 112.98 -6.76 112.99 ;
      RECT  -12.79 113.32 -12.45 113.64 ;
      RECT  -7.09 113.19 -6.76 113.31 ;
      RECT  -2.31 114.35 -1.78 114.58 ;
      RECT  -14.53 110.34 -1.4 110.75 ;
      RECT  -13.41 112.09 -11.96 112.29 ;
      RECT  -12.25 112.99 -6.76 113.19 ;
      RECT  -12.9 110.75 -12.49 111.12 ;
      RECT  -10.75 110.75 -10.34 111.12 ;
      RECT  -11.17 112.49 -6.25 112.74 ;
      RECT  -11.7 112.29 -11.4 112.35 ;
      RECT  -3.66 114.35 -3.13 114.58 ;
      RECT  -5.43 114.35 -4.9 114.58 ;
      RECT  -4.95 110.75 -4.54 111.12 ;
      RECT  -5.37 112.98 -5.04 112.99 ;
      RECT  -5.37 113.19 -5.04 113.31 ;
      RECT  -5.9 112.09 -2.23 112.29 ;
      RECT  -13.41 112.29 -13.12 112.35 ;
      RECT  -11.86 110.75 -11.45 111.12 ;
      RECT  -5.9 112.29 -5.6 112.33 ;
      RECT  -6.45 112.99 -5.04 113.19 ;
      RECT  -8.6 111.98 -8.27 112.08 ;
      RECT  -11.17 112.74 -10.84 112.77 ;
      RECT  -2.57 111.99 -2.23 112.09 ;
      RECT  -6.06 110.75 -5.65 111.12 ;
      RECT  -4.23 112.64 -3.6 112.96 ;
      RECT  -11.23 114.35 -10.7 114.58 ;
      RECT  -6.49 112.0 -6.16 112.33 ;
      RECT  -11.17 112.44 -10.84 112.49 ;
      RECT  -3.85 110.75 -3.44 111.12 ;
      RECT  -11.7 112.08 -8.27 112.29 ;
      RECT  -11.7 112.04 -11.4 112.08 ;
      RECT  -2.57 112.29 -2.23 112.32 ;
      RECT  -12.75 114.35 -12.22 114.58 ;
      RECT  -12.29 112.04 -11.96 112.09 ;
      RECT  -7.1 110.75 -6.69 111.12 ;
      RECT  -6.45 112.74 -6.25 112.99 ;
      RECT  -13.41 112.06 -13.12 112.09 ;
      RECT  -5.9 112.02 -5.6 112.09 ;
      RECT  -6.95 115.25 -6.42 115.02 ;
      RECT  -11.17 116.41 -10.84 116.29 ;
      RECT  -6.45 117.27 -6.25 117.11 ;
      RECT  -8.6 117.31 -8.27 117.29 ;
      RECT  -14.28 117.52 -13.97 117.2 ;
      RECT  -14.53 115.02 -1.4 114.57 ;
      RECT  -12.29 117.31 -11.96 117.23 ;
      RECT  -11.17 116.62 -10.84 116.61 ;
      RECT  -12.25 117.23 -12.05 116.61 ;
      RECT  -9.71 115.25 -9.18 115.02 ;
      RECT  -7.09 116.62 -6.76 116.61 ;
      RECT  -12.79 116.28 -12.45 115.96 ;
      RECT  -7.09 116.41 -6.76 116.29 ;
      RECT  -2.31 115.25 -1.78 115.02 ;
      RECT  -14.53 119.26 -1.4 118.85 ;
      RECT  -13.41 117.51 -11.96 117.31 ;
      RECT  -12.25 116.61 -6.76 116.41 ;
      RECT  -12.9 118.85 -12.49 118.48 ;
      RECT  -10.75 118.85 -10.34 118.48 ;
      RECT  -11.17 117.11 -6.25 116.86 ;
      RECT  -11.7 117.31 -11.4 117.25 ;
      RECT  -3.66 115.25 -3.13 115.02 ;
      RECT  -5.43 115.25 -4.9 115.02 ;
      RECT  -4.95 118.85 -4.54 118.48 ;
      RECT  -5.37 116.62 -5.04 116.61 ;
      RECT  -5.37 116.41 -5.04 116.29 ;
      RECT  -5.9 117.51 -2.23 117.31 ;
      RECT  -13.41 117.31 -13.12 117.25 ;
      RECT  -11.86 118.85 -11.45 118.48 ;
      RECT  -5.9 117.31 -5.6 117.27 ;
      RECT  -6.45 116.61 -5.04 116.41 ;
      RECT  -8.6 117.62 -8.27 117.52 ;
      RECT  -11.17 116.86 -10.84 116.83 ;
      RECT  -2.57 117.61 -2.23 117.51 ;
      RECT  -6.06 118.85 -5.65 118.48 ;
      RECT  -4.23 116.96 -3.6 116.64 ;
      RECT  -11.23 115.25 -10.7 115.02 ;
      RECT  -6.49 117.6 -6.16 117.27 ;
      RECT  -11.17 117.16 -10.84 117.11 ;
      RECT  -3.85 118.85 -3.44 118.48 ;
      RECT  -11.7 117.52 -8.27 117.31 ;
      RECT  -11.7 117.56 -11.4 117.52 ;
      RECT  -2.57 117.31 -2.23 117.28 ;
      RECT  -12.75 115.25 -12.22 115.02 ;
      RECT  -12.29 117.56 -11.96 117.51 ;
      RECT  -7.1 118.85 -6.69 118.48 ;
      RECT  -6.45 116.86 -6.25 116.61 ;
      RECT  -13.41 117.54 -13.12 117.51 ;
      RECT  -5.9 117.58 -5.6 117.51 ;
      RECT  19.31 -6.25 19.84 -6.02 ;
      RECT  15.09 -7.41 15.42 -7.29 ;
      RECT  19.81 -8.27 20.01 -8.11 ;
      RECT  17.66 -8.31 17.99 -8.29 ;
      RECT  11.98 -8.52 12.29 -8.2 ;
      RECT  11.73 -6.02 24.86 -5.57 ;
      RECT  13.97 -8.31 14.3 -8.23 ;
      RECT  15.09 -7.62 15.42 -7.61 ;
      RECT  14.01 -8.23 14.21 -7.61 ;
      RECT  16.55 -6.25 17.08 -6.02 ;
      RECT  19.17 -7.62 19.5 -7.61 ;
      RECT  13.47 -7.28 13.81 -6.96 ;
      RECT  19.17 -7.41 19.5 -7.29 ;
      RECT  23.95 -6.25 24.48 -6.02 ;
      RECT  11.73 -10.26 24.86 -9.85 ;
      RECT  12.85 -8.51 14.3 -8.31 ;
      RECT  14.01 -7.61 19.5 -7.41 ;
      RECT  13.36 -9.85 13.77 -9.48 ;
      RECT  15.51 -9.85 15.92 -9.48 ;
      RECT  15.09 -8.11 20.01 -7.86 ;
      RECT  14.56 -8.31 14.86 -8.25 ;
      RECT  22.6 -6.25 23.13 -6.02 ;
      RECT  20.83 -6.25 21.36 -6.02 ;
      RECT  21.31 -9.85 21.72 -9.48 ;
      RECT  20.89 -7.62 21.22 -7.61 ;
      RECT  20.89 -7.41 21.22 -7.29 ;
      RECT  20.36 -8.51 24.03 -8.31 ;
      RECT  12.85 -8.31 13.14 -8.25 ;
      RECT  14.4 -9.85 14.81 -9.48 ;
      RECT  20.36 -8.31 20.66 -8.27 ;
      RECT  19.81 -7.61 21.22 -7.41 ;
      RECT  17.66 -8.62 17.99 -8.52 ;
      RECT  15.09 -7.86 15.42 -7.83 ;
      RECT  23.69 -8.61 24.03 -8.51 ;
      RECT  20.2 -9.85 20.61 -9.48 ;
      RECT  22.03 -7.96 22.66 -7.64 ;
      RECT  15.03 -6.25 15.56 -6.02 ;
      RECT  19.77 -8.6 20.1 -8.27 ;
      RECT  15.09 -8.16 15.42 -8.11 ;
      RECT  22.41 -9.85 22.82 -9.48 ;
      RECT  14.56 -8.52 17.99 -8.31 ;
      RECT  14.56 -8.56 14.86 -8.52 ;
      RECT  23.69 -8.31 24.03 -8.28 ;
      RECT  13.51 -6.25 14.04 -6.02 ;
      RECT  13.97 -8.56 14.3 -8.51 ;
      RECT  19.16 -9.85 19.57 -9.48 ;
      RECT  19.81 -7.86 20.01 -7.61 ;
      RECT  12.85 -8.54 13.14 -8.51 ;
      RECT  20.36 -8.58 20.66 -8.51 ;
      RECT  32.44 -6.25 32.97 -6.02 ;
      RECT  28.22 -7.41 28.55 -7.29 ;
      RECT  32.94 -8.27 33.14 -8.11 ;
      RECT  30.79 -8.31 31.12 -8.29 ;
      RECT  25.11 -8.52 25.42 -8.2 ;
      RECT  24.86 -6.02 37.99 -5.57 ;
      RECT  27.1 -8.31 27.43 -8.23 ;
      RECT  28.22 -7.62 28.55 -7.61 ;
      RECT  27.14 -8.23 27.34 -7.61 ;
      RECT  29.68 -6.25 30.21 -6.02 ;
      RECT  32.3 -7.62 32.63 -7.61 ;
      RECT  26.6 -7.28 26.94 -6.96 ;
      RECT  32.3 -7.41 32.63 -7.29 ;
      RECT  37.08 -6.25 37.61 -6.02 ;
      RECT  24.86 -10.26 37.99 -9.85 ;
      RECT  25.98 -8.51 27.43 -8.31 ;
      RECT  27.14 -7.61 32.63 -7.41 ;
      RECT  26.49 -9.85 26.9 -9.48 ;
      RECT  28.64 -9.85 29.05 -9.48 ;
      RECT  28.22 -8.11 33.14 -7.86 ;
      RECT  27.69 -8.31 27.99 -8.25 ;
      RECT  35.73 -6.25 36.26 -6.02 ;
      RECT  33.96 -6.25 34.49 -6.02 ;
      RECT  34.44 -9.85 34.85 -9.48 ;
      RECT  34.02 -7.62 34.35 -7.61 ;
      RECT  34.02 -7.41 34.35 -7.29 ;
      RECT  33.49 -8.51 37.16 -8.31 ;
      RECT  25.98 -8.31 26.27 -8.25 ;
      RECT  27.53 -9.85 27.94 -9.48 ;
      RECT  33.49 -8.31 33.79 -8.27 ;
      RECT  32.94 -7.61 34.35 -7.41 ;
      RECT  30.79 -8.62 31.12 -8.52 ;
      RECT  28.22 -7.86 28.55 -7.83 ;
      RECT  36.82 -8.61 37.16 -8.51 ;
      RECT  33.33 -9.85 33.74 -9.48 ;
      RECT  35.16 -7.96 35.79 -7.64 ;
      RECT  28.16 -6.25 28.69 -6.02 ;
      RECT  32.9 -8.6 33.23 -8.27 ;
      RECT  28.22 -8.16 28.55 -8.11 ;
      RECT  35.54 -9.85 35.95 -9.48 ;
      RECT  27.69 -8.52 31.12 -8.31 ;
      RECT  27.69 -8.56 27.99 -8.52 ;
      RECT  36.82 -8.31 37.16 -8.28 ;
      RECT  26.64 -6.25 27.17 -6.02 ;
      RECT  27.1 -8.56 27.43 -8.51 ;
      RECT  32.29 -9.85 32.7 -9.48 ;
      RECT  32.94 -7.86 33.14 -7.61 ;
      RECT  25.98 -8.54 26.27 -8.51 ;
      RECT  33.49 -8.58 33.79 -8.51 ;
   LAYER  m2 ;
      RECT  56.45 36.51 56.77 36.62 ;
      RECT  56.96 36.52 57.28 36.62 ;
      RECT  56.45 36.3 56.77 36.37 ;
      RECT  56.96 36.3 57.28 36.38 ;
      RECT  56.12 35.66 56.26 36.37 ;
      RECT  56.12 36.37 56.77 36.51 ;
      RECT  56.96 36.38 57.68 36.52 ;
      RECT  56.12 36.51 56.26 41.4 ;
      RECT  57.54 35.66 57.68 36.38 ;
      RECT  57.54 36.52 57.68 41.4 ;
      RECT  56.45 45.85 56.77 45.74 ;
      RECT  56.96 45.84 57.28 45.74 ;
      RECT  56.45 46.06 56.77 45.99 ;
      RECT  56.96 46.06 57.28 45.98 ;
      RECT  56.12 46.7 56.26 45.99 ;
      RECT  56.12 45.99 56.77 45.85 ;
      RECT  56.96 45.98 57.68 45.84 ;
      RECT  56.12 45.85 56.26 40.96 ;
      RECT  57.54 46.7 57.68 45.98 ;
      RECT  57.54 45.84 57.68 40.96 ;
      RECT  56.45 47.15 56.77 47.26 ;
      RECT  56.96 47.16 57.28 47.26 ;
      RECT  56.45 46.94 56.77 47.01 ;
      RECT  56.96 46.94 57.28 47.02 ;
      RECT  56.12 46.3 56.26 47.01 ;
      RECT  56.12 47.01 56.77 47.15 ;
      RECT  56.96 47.02 57.68 47.16 ;
      RECT  56.12 47.15 56.26 52.04 ;
      RECT  57.54 46.3 57.68 47.02 ;
      RECT  57.54 47.16 57.68 52.04 ;
      RECT  56.45 56.49 56.77 56.38 ;
      RECT  56.96 56.48 57.28 56.38 ;
      RECT  56.45 56.7 56.77 56.63 ;
      RECT  56.96 56.7 57.28 56.62 ;
      RECT  56.12 57.34 56.26 56.63 ;
      RECT  56.12 56.63 56.77 56.49 ;
      RECT  56.96 56.62 57.68 56.48 ;
      RECT  56.12 56.49 56.26 51.6 ;
      RECT  57.54 57.34 57.68 56.62 ;
      RECT  57.54 56.48 57.68 51.6 ;
      RECT  56.45 57.79 56.77 57.9 ;
      RECT  56.96 57.8 57.28 57.9 ;
      RECT  56.45 57.58 56.77 57.65 ;
      RECT  56.96 57.58 57.28 57.66 ;
      RECT  56.12 56.94 56.26 57.65 ;
      RECT  56.12 57.65 56.77 57.79 ;
      RECT  56.96 57.66 57.68 57.8 ;
      RECT  56.12 57.79 56.26 62.68 ;
      RECT  57.54 56.94 57.68 57.66 ;
      RECT  57.54 57.8 57.68 62.68 ;
      RECT  56.45 67.13 56.77 67.02 ;
      RECT  56.96 67.12 57.28 67.02 ;
      RECT  56.45 67.34 56.77 67.27 ;
      RECT  56.96 67.34 57.28 67.26 ;
      RECT  56.12 67.98 56.26 67.27 ;
      RECT  56.12 67.27 56.77 67.13 ;
      RECT  56.96 67.26 57.68 67.12 ;
      RECT  56.12 67.13 56.26 62.24 ;
      RECT  57.54 67.98 57.68 67.26 ;
      RECT  57.54 67.12 57.68 62.24 ;
      RECT  56.45 68.43 56.77 68.54 ;
      RECT  56.96 68.44 57.28 68.54 ;
      RECT  56.45 68.22 56.77 68.29 ;
      RECT  56.96 68.22 57.28 68.3 ;
      RECT  56.12 67.58 56.26 68.29 ;
      RECT  56.12 68.29 56.77 68.43 ;
      RECT  56.96 68.3 57.68 68.44 ;
      RECT  56.12 68.43 56.26 73.32 ;
      RECT  57.54 67.58 57.68 68.3 ;
      RECT  57.54 68.44 57.68 73.32 ;
      RECT  56.45 77.77 56.77 77.66 ;
      RECT  56.96 77.76 57.28 77.66 ;
      RECT  56.45 77.98 56.77 77.91 ;
      RECT  56.96 77.98 57.28 77.9 ;
      RECT  56.12 78.62 56.26 77.91 ;
      RECT  56.12 77.91 56.77 77.77 ;
      RECT  56.96 77.9 57.68 77.76 ;
      RECT  56.12 77.77 56.26 72.88 ;
      RECT  57.54 78.62 57.68 77.9 ;
      RECT  57.54 77.76 57.68 72.88 ;
      RECT  56.45 79.07 56.77 79.18 ;
      RECT  56.96 79.08 57.28 79.18 ;
      RECT  56.45 78.86 56.77 78.93 ;
      RECT  56.96 78.86 57.28 78.94 ;
      RECT  56.12 78.22 56.26 78.93 ;
      RECT  56.12 78.93 56.77 79.07 ;
      RECT  56.96 78.94 57.68 79.08 ;
      RECT  56.12 79.07 56.26 83.96 ;
      RECT  57.54 78.22 57.68 78.94 ;
      RECT  57.54 79.08 57.68 83.96 ;
      RECT  56.45 88.41 56.77 88.3 ;
      RECT  56.96 88.4 57.28 88.3 ;
      RECT  56.45 88.62 56.77 88.55 ;
      RECT  56.96 88.62 57.28 88.54 ;
      RECT  56.12 89.26 56.26 88.55 ;
      RECT  56.12 88.55 56.77 88.41 ;
      RECT  56.96 88.54 57.68 88.4 ;
      RECT  56.12 88.41 56.26 83.52 ;
      RECT  57.54 89.26 57.68 88.54 ;
      RECT  57.54 88.4 57.68 83.52 ;
      RECT  56.45 89.71 56.77 89.82 ;
      RECT  56.96 89.72 57.28 89.82 ;
      RECT  56.45 89.5 56.77 89.57 ;
      RECT  56.96 89.5 57.28 89.58 ;
      RECT  56.12 88.86 56.26 89.57 ;
      RECT  56.12 89.57 56.77 89.71 ;
      RECT  56.96 89.58 57.68 89.72 ;
      RECT  56.12 89.71 56.26 94.6 ;
      RECT  57.54 88.86 57.68 89.58 ;
      RECT  57.54 89.72 57.68 94.6 ;
      RECT  56.45 99.05 56.77 98.94 ;
      RECT  56.96 99.04 57.28 98.94 ;
      RECT  56.45 99.26 56.77 99.19 ;
      RECT  56.96 99.26 57.28 99.18 ;
      RECT  56.12 99.9 56.26 99.19 ;
      RECT  56.12 99.19 56.77 99.05 ;
      RECT  56.96 99.18 57.68 99.04 ;
      RECT  56.12 99.05 56.26 94.16 ;
      RECT  57.54 99.9 57.68 99.18 ;
      RECT  57.54 99.04 57.68 94.16 ;
      RECT  56.45 100.35 56.77 100.46 ;
      RECT  56.96 100.36 57.28 100.46 ;
      RECT  56.45 100.14 56.77 100.21 ;
      RECT  56.96 100.14 57.28 100.22 ;
      RECT  56.12 99.5 56.26 100.21 ;
      RECT  56.12 100.21 56.77 100.35 ;
      RECT  56.96 100.22 57.68 100.36 ;
      RECT  56.12 100.35 56.26 105.24 ;
      RECT  57.54 99.5 57.68 100.22 ;
      RECT  57.54 100.36 57.68 105.24 ;
      RECT  56.45 109.69 56.77 109.58 ;
      RECT  56.96 109.68 57.28 109.58 ;
      RECT  56.45 109.9 56.77 109.83 ;
      RECT  56.96 109.9 57.28 109.82 ;
      RECT  56.12 110.54 56.26 109.83 ;
      RECT  56.12 109.83 56.77 109.69 ;
      RECT  56.96 109.82 57.68 109.68 ;
      RECT  56.12 109.69 56.26 104.8 ;
      RECT  57.54 110.54 57.68 109.82 ;
      RECT  57.54 109.68 57.68 104.8 ;
      RECT  56.45 110.99 56.77 111.1 ;
      RECT  56.96 111.0 57.28 111.1 ;
      RECT  56.45 110.78 56.77 110.85 ;
      RECT  56.96 110.78 57.28 110.86 ;
      RECT  56.12 110.14 56.26 110.85 ;
      RECT  56.12 110.85 56.77 110.99 ;
      RECT  56.96 110.86 57.68 111.0 ;
      RECT  56.12 110.99 56.26 115.88 ;
      RECT  57.54 110.14 57.68 110.86 ;
      RECT  57.54 111.0 57.68 115.88 ;
      RECT  56.45 120.33 56.77 120.22 ;
      RECT  56.96 120.32 57.28 120.22 ;
      RECT  56.45 120.54 56.77 120.47 ;
      RECT  56.96 120.54 57.28 120.46 ;
      RECT  56.12 121.18 56.26 120.47 ;
      RECT  56.12 120.47 56.77 120.33 ;
      RECT  56.96 120.46 57.68 120.32 ;
      RECT  56.12 120.33 56.26 115.44 ;
      RECT  57.54 121.18 57.68 120.46 ;
      RECT  57.54 120.32 57.68 115.44 ;
      RECT  60.45 36.51 60.77 36.62 ;
      RECT  60.96 36.52 61.28 36.62 ;
      RECT  60.45 36.3 60.77 36.37 ;
      RECT  60.96 36.3 61.28 36.38 ;
      RECT  60.12 35.66 60.26 36.37 ;
      RECT  60.12 36.37 60.77 36.51 ;
      RECT  60.96 36.38 61.68 36.52 ;
      RECT  60.12 36.51 60.26 41.4 ;
      RECT  61.54 35.66 61.68 36.38 ;
      RECT  61.54 36.52 61.68 41.4 ;
      RECT  60.45 45.85 60.77 45.74 ;
      RECT  60.96 45.84 61.28 45.74 ;
      RECT  60.45 46.06 60.77 45.99 ;
      RECT  60.96 46.06 61.28 45.98 ;
      RECT  60.12 46.7 60.26 45.99 ;
      RECT  60.12 45.99 60.77 45.85 ;
      RECT  60.96 45.98 61.68 45.84 ;
      RECT  60.12 45.85 60.26 40.96 ;
      RECT  61.54 46.7 61.68 45.98 ;
      RECT  61.54 45.84 61.68 40.96 ;
      RECT  60.45 47.15 60.77 47.26 ;
      RECT  60.96 47.16 61.28 47.26 ;
      RECT  60.45 46.94 60.77 47.01 ;
      RECT  60.96 46.94 61.28 47.02 ;
      RECT  60.12 46.3 60.26 47.01 ;
      RECT  60.12 47.01 60.77 47.15 ;
      RECT  60.96 47.02 61.68 47.16 ;
      RECT  60.12 47.15 60.26 52.04 ;
      RECT  61.54 46.3 61.68 47.02 ;
      RECT  61.54 47.16 61.68 52.04 ;
      RECT  60.45 56.49 60.77 56.38 ;
      RECT  60.96 56.48 61.28 56.38 ;
      RECT  60.45 56.7 60.77 56.63 ;
      RECT  60.96 56.7 61.28 56.62 ;
      RECT  60.12 57.34 60.26 56.63 ;
      RECT  60.12 56.63 60.77 56.49 ;
      RECT  60.96 56.62 61.68 56.48 ;
      RECT  60.12 56.49 60.26 51.6 ;
      RECT  61.54 57.34 61.68 56.62 ;
      RECT  61.54 56.48 61.68 51.6 ;
      RECT  60.45 57.79 60.77 57.9 ;
      RECT  60.96 57.8 61.28 57.9 ;
      RECT  60.45 57.58 60.77 57.65 ;
      RECT  60.96 57.58 61.28 57.66 ;
      RECT  60.12 56.94 60.26 57.65 ;
      RECT  60.12 57.65 60.77 57.79 ;
      RECT  60.96 57.66 61.68 57.8 ;
      RECT  60.12 57.79 60.26 62.68 ;
      RECT  61.54 56.94 61.68 57.66 ;
      RECT  61.54 57.8 61.68 62.68 ;
      RECT  60.45 67.13 60.77 67.02 ;
      RECT  60.96 67.12 61.28 67.02 ;
      RECT  60.45 67.34 60.77 67.27 ;
      RECT  60.96 67.34 61.28 67.26 ;
      RECT  60.12 67.98 60.26 67.27 ;
      RECT  60.12 67.27 60.77 67.13 ;
      RECT  60.96 67.26 61.68 67.12 ;
      RECT  60.12 67.13 60.26 62.24 ;
      RECT  61.54 67.98 61.68 67.26 ;
      RECT  61.54 67.12 61.68 62.24 ;
      RECT  60.45 68.43 60.77 68.54 ;
      RECT  60.96 68.44 61.28 68.54 ;
      RECT  60.45 68.22 60.77 68.29 ;
      RECT  60.96 68.22 61.28 68.3 ;
      RECT  60.12 67.58 60.26 68.29 ;
      RECT  60.12 68.29 60.77 68.43 ;
      RECT  60.96 68.3 61.68 68.44 ;
      RECT  60.12 68.43 60.26 73.32 ;
      RECT  61.54 67.58 61.68 68.3 ;
      RECT  61.54 68.44 61.68 73.32 ;
      RECT  60.45 77.77 60.77 77.66 ;
      RECT  60.96 77.76 61.28 77.66 ;
      RECT  60.45 77.98 60.77 77.91 ;
      RECT  60.96 77.98 61.28 77.9 ;
      RECT  60.12 78.62 60.26 77.91 ;
      RECT  60.12 77.91 60.77 77.77 ;
      RECT  60.96 77.9 61.68 77.76 ;
      RECT  60.12 77.77 60.26 72.88 ;
      RECT  61.54 78.62 61.68 77.9 ;
      RECT  61.54 77.76 61.68 72.88 ;
      RECT  60.45 79.07 60.77 79.18 ;
      RECT  60.96 79.08 61.28 79.18 ;
      RECT  60.45 78.86 60.77 78.93 ;
      RECT  60.96 78.86 61.28 78.94 ;
      RECT  60.12 78.22 60.26 78.93 ;
      RECT  60.12 78.93 60.77 79.07 ;
      RECT  60.96 78.94 61.68 79.08 ;
      RECT  60.12 79.07 60.26 83.96 ;
      RECT  61.54 78.22 61.68 78.94 ;
      RECT  61.54 79.08 61.68 83.96 ;
      RECT  60.45 88.41 60.77 88.3 ;
      RECT  60.96 88.4 61.28 88.3 ;
      RECT  60.45 88.62 60.77 88.55 ;
      RECT  60.96 88.62 61.28 88.54 ;
      RECT  60.12 89.26 60.26 88.55 ;
      RECT  60.12 88.55 60.77 88.41 ;
      RECT  60.96 88.54 61.68 88.4 ;
      RECT  60.12 88.41 60.26 83.52 ;
      RECT  61.54 89.26 61.68 88.54 ;
      RECT  61.54 88.4 61.68 83.52 ;
      RECT  60.45 89.71 60.77 89.82 ;
      RECT  60.96 89.72 61.28 89.82 ;
      RECT  60.45 89.5 60.77 89.57 ;
      RECT  60.96 89.5 61.28 89.58 ;
      RECT  60.12 88.86 60.26 89.57 ;
      RECT  60.12 89.57 60.77 89.71 ;
      RECT  60.96 89.58 61.68 89.72 ;
      RECT  60.12 89.71 60.26 94.6 ;
      RECT  61.54 88.86 61.68 89.58 ;
      RECT  61.54 89.72 61.68 94.6 ;
      RECT  60.45 99.05 60.77 98.94 ;
      RECT  60.96 99.04 61.28 98.94 ;
      RECT  60.45 99.26 60.77 99.19 ;
      RECT  60.96 99.26 61.28 99.18 ;
      RECT  60.12 99.9 60.26 99.19 ;
      RECT  60.12 99.19 60.77 99.05 ;
      RECT  60.96 99.18 61.68 99.04 ;
      RECT  60.12 99.05 60.26 94.16 ;
      RECT  61.54 99.9 61.68 99.18 ;
      RECT  61.54 99.04 61.68 94.16 ;
      RECT  60.45 100.35 60.77 100.46 ;
      RECT  60.96 100.36 61.28 100.46 ;
      RECT  60.45 100.14 60.77 100.21 ;
      RECT  60.96 100.14 61.28 100.22 ;
      RECT  60.12 99.5 60.26 100.21 ;
      RECT  60.12 100.21 60.77 100.35 ;
      RECT  60.96 100.22 61.68 100.36 ;
      RECT  60.12 100.35 60.26 105.24 ;
      RECT  61.54 99.5 61.68 100.22 ;
      RECT  61.54 100.36 61.68 105.24 ;
      RECT  60.45 109.69 60.77 109.58 ;
      RECT  60.96 109.68 61.28 109.58 ;
      RECT  60.45 109.9 60.77 109.83 ;
      RECT  60.96 109.9 61.28 109.82 ;
      RECT  60.12 110.54 60.26 109.83 ;
      RECT  60.12 109.83 60.77 109.69 ;
      RECT  60.96 109.82 61.68 109.68 ;
      RECT  60.12 109.69 60.26 104.8 ;
      RECT  61.54 110.54 61.68 109.82 ;
      RECT  61.54 109.68 61.68 104.8 ;
      RECT  60.45 110.99 60.77 111.1 ;
      RECT  60.96 111.0 61.28 111.1 ;
      RECT  60.45 110.78 60.77 110.85 ;
      RECT  60.96 110.78 61.28 110.86 ;
      RECT  60.12 110.14 60.26 110.85 ;
      RECT  60.12 110.85 60.77 110.99 ;
      RECT  60.96 110.86 61.68 111.0 ;
      RECT  60.12 110.99 60.26 115.88 ;
      RECT  61.54 110.14 61.68 110.86 ;
      RECT  61.54 111.0 61.68 115.88 ;
      RECT  60.45 120.33 60.77 120.22 ;
      RECT  60.96 120.32 61.28 120.22 ;
      RECT  60.45 120.54 60.77 120.47 ;
      RECT  60.96 120.54 61.28 120.46 ;
      RECT  60.12 121.18 60.26 120.47 ;
      RECT  60.12 120.47 60.77 120.33 ;
      RECT  60.96 120.46 61.68 120.32 ;
      RECT  60.12 120.33 60.26 115.44 ;
      RECT  61.54 121.18 61.68 120.46 ;
      RECT  61.54 120.32 61.68 115.44 ;
      RECT  56.12 35.86 56.77 120.98 ;
      RECT  56.96 35.86 57.68 120.98 ;
      RECT  60.12 35.86 60.77 120.98 ;
      RECT  60.96 35.86 61.68 120.98 ;
      RECT  52.12 25.02 52.26 30.76 ;
      RECT  53.54 25.02 53.68 30.76 ;
      RECT  52.45 35.21 52.77 35.1 ;
      RECT  52.96 35.2 53.28 35.1 ;
      RECT  52.45 35.42 52.77 35.35 ;
      RECT  52.96 35.42 53.28 35.34 ;
      RECT  52.12 36.06 52.26 35.35 ;
      RECT  52.12 35.35 52.77 35.21 ;
      RECT  52.96 35.34 53.68 35.2 ;
      RECT  52.12 35.21 52.26 30.32 ;
      RECT  53.54 36.06 53.68 35.34 ;
      RECT  53.54 35.2 53.68 30.32 ;
      RECT  52.45 36.51 52.77 36.62 ;
      RECT  52.96 36.52 53.28 36.62 ;
      RECT  52.45 36.3 52.77 36.37 ;
      RECT  52.96 36.3 53.28 36.38 ;
      RECT  52.12 35.66 52.26 36.37 ;
      RECT  52.12 36.37 52.77 36.51 ;
      RECT  52.96 36.38 53.68 36.52 ;
      RECT  52.12 36.51 52.26 41.4 ;
      RECT  53.54 35.66 53.68 36.38 ;
      RECT  53.54 36.52 53.68 41.4 ;
      RECT  52.45 45.85 52.77 45.74 ;
      RECT  52.96 45.84 53.28 45.74 ;
      RECT  52.45 46.06 52.77 45.99 ;
      RECT  52.96 46.06 53.28 45.98 ;
      RECT  52.12 46.7 52.26 45.99 ;
      RECT  52.12 45.99 52.77 45.85 ;
      RECT  52.96 45.98 53.68 45.84 ;
      RECT  52.12 45.85 52.26 40.96 ;
      RECT  53.54 46.7 53.68 45.98 ;
      RECT  53.54 45.84 53.68 40.96 ;
      RECT  52.45 47.15 52.77 47.26 ;
      RECT  52.96 47.16 53.28 47.26 ;
      RECT  52.45 46.94 52.77 47.01 ;
      RECT  52.96 46.94 53.28 47.02 ;
      RECT  52.12 46.3 52.26 47.01 ;
      RECT  52.12 47.01 52.77 47.15 ;
      RECT  52.96 47.02 53.68 47.16 ;
      RECT  52.12 47.15 52.26 52.04 ;
      RECT  53.54 46.3 53.68 47.02 ;
      RECT  53.54 47.16 53.68 52.04 ;
      RECT  52.45 56.49 52.77 56.38 ;
      RECT  52.96 56.48 53.28 56.38 ;
      RECT  52.45 56.7 52.77 56.63 ;
      RECT  52.96 56.7 53.28 56.62 ;
      RECT  52.12 57.34 52.26 56.63 ;
      RECT  52.12 56.63 52.77 56.49 ;
      RECT  52.96 56.62 53.68 56.48 ;
      RECT  52.12 56.49 52.26 51.6 ;
      RECT  53.54 57.34 53.68 56.62 ;
      RECT  53.54 56.48 53.68 51.6 ;
      RECT  52.45 57.79 52.77 57.9 ;
      RECT  52.96 57.8 53.28 57.9 ;
      RECT  52.45 57.58 52.77 57.65 ;
      RECT  52.96 57.58 53.28 57.66 ;
      RECT  52.12 56.94 52.26 57.65 ;
      RECT  52.12 57.65 52.77 57.79 ;
      RECT  52.96 57.66 53.68 57.8 ;
      RECT  52.12 57.79 52.26 62.68 ;
      RECT  53.54 56.94 53.68 57.66 ;
      RECT  53.54 57.8 53.68 62.68 ;
      RECT  52.45 67.13 52.77 67.02 ;
      RECT  52.96 67.12 53.28 67.02 ;
      RECT  52.45 67.34 52.77 67.27 ;
      RECT  52.96 67.34 53.28 67.26 ;
      RECT  52.12 67.98 52.26 67.27 ;
      RECT  52.12 67.27 52.77 67.13 ;
      RECT  52.96 67.26 53.68 67.12 ;
      RECT  52.12 67.13 52.26 62.24 ;
      RECT  53.54 67.98 53.68 67.26 ;
      RECT  53.54 67.12 53.68 62.24 ;
      RECT  52.45 68.43 52.77 68.54 ;
      RECT  52.96 68.44 53.28 68.54 ;
      RECT  52.45 68.22 52.77 68.29 ;
      RECT  52.96 68.22 53.28 68.3 ;
      RECT  52.12 67.58 52.26 68.29 ;
      RECT  52.12 68.29 52.77 68.43 ;
      RECT  52.96 68.3 53.68 68.44 ;
      RECT  52.12 68.43 52.26 73.32 ;
      RECT  53.54 67.58 53.68 68.3 ;
      RECT  53.54 68.44 53.68 73.32 ;
      RECT  52.45 77.77 52.77 77.66 ;
      RECT  52.96 77.76 53.28 77.66 ;
      RECT  52.45 77.98 52.77 77.91 ;
      RECT  52.96 77.98 53.28 77.9 ;
      RECT  52.12 78.62 52.26 77.91 ;
      RECT  52.12 77.91 52.77 77.77 ;
      RECT  52.96 77.9 53.68 77.76 ;
      RECT  52.12 77.77 52.26 72.88 ;
      RECT  53.54 78.62 53.68 77.9 ;
      RECT  53.54 77.76 53.68 72.88 ;
      RECT  52.45 79.07 52.77 79.18 ;
      RECT  52.96 79.08 53.28 79.18 ;
      RECT  52.45 78.86 52.77 78.93 ;
      RECT  52.96 78.86 53.28 78.94 ;
      RECT  52.12 78.22 52.26 78.93 ;
      RECT  52.12 78.93 52.77 79.07 ;
      RECT  52.96 78.94 53.68 79.08 ;
      RECT  52.12 79.07 52.26 83.96 ;
      RECT  53.54 78.22 53.68 78.94 ;
      RECT  53.54 79.08 53.68 83.96 ;
      RECT  52.45 88.41 52.77 88.3 ;
      RECT  52.96 88.4 53.28 88.3 ;
      RECT  52.45 88.62 52.77 88.55 ;
      RECT  52.96 88.62 53.28 88.54 ;
      RECT  52.12 89.26 52.26 88.55 ;
      RECT  52.12 88.55 52.77 88.41 ;
      RECT  52.96 88.54 53.68 88.4 ;
      RECT  52.12 88.41 52.26 83.52 ;
      RECT  53.54 89.26 53.68 88.54 ;
      RECT  53.54 88.4 53.68 83.52 ;
      RECT  52.45 89.71 52.77 89.82 ;
      RECT  52.96 89.72 53.28 89.82 ;
      RECT  52.45 89.5 52.77 89.57 ;
      RECT  52.96 89.5 53.28 89.58 ;
      RECT  52.12 88.86 52.26 89.57 ;
      RECT  52.12 89.57 52.77 89.71 ;
      RECT  52.96 89.58 53.68 89.72 ;
      RECT  52.12 89.71 52.26 94.6 ;
      RECT  53.54 88.86 53.68 89.58 ;
      RECT  53.54 89.72 53.68 94.6 ;
      RECT  52.45 99.05 52.77 98.94 ;
      RECT  52.96 99.04 53.28 98.94 ;
      RECT  52.45 99.26 52.77 99.19 ;
      RECT  52.96 99.26 53.28 99.18 ;
      RECT  52.12 99.9 52.26 99.19 ;
      RECT  52.12 99.19 52.77 99.05 ;
      RECT  52.96 99.18 53.68 99.04 ;
      RECT  52.12 99.05 52.26 94.16 ;
      RECT  53.54 99.9 53.68 99.18 ;
      RECT  53.54 99.04 53.68 94.16 ;
      RECT  52.45 100.35 52.77 100.46 ;
      RECT  52.96 100.36 53.28 100.46 ;
      RECT  52.45 100.14 52.77 100.21 ;
      RECT  52.96 100.14 53.28 100.22 ;
      RECT  52.12 99.5 52.26 100.21 ;
      RECT  52.12 100.21 52.77 100.35 ;
      RECT  52.96 100.22 53.68 100.36 ;
      RECT  52.12 100.35 52.26 105.24 ;
      RECT  53.54 99.5 53.68 100.22 ;
      RECT  53.54 100.36 53.68 105.24 ;
      RECT  52.45 109.69 52.77 109.58 ;
      RECT  52.96 109.68 53.28 109.58 ;
      RECT  52.45 109.9 52.77 109.83 ;
      RECT  52.96 109.9 53.28 109.82 ;
      RECT  52.12 110.54 52.26 109.83 ;
      RECT  52.12 109.83 52.77 109.69 ;
      RECT  52.96 109.82 53.68 109.68 ;
      RECT  52.12 109.69 52.26 104.8 ;
      RECT  53.54 110.54 53.68 109.82 ;
      RECT  53.54 109.68 53.68 104.8 ;
      RECT  52.45 110.99 52.77 111.1 ;
      RECT  52.96 111.0 53.28 111.1 ;
      RECT  52.45 110.78 52.77 110.85 ;
      RECT  52.96 110.78 53.28 110.86 ;
      RECT  52.12 110.14 52.26 110.85 ;
      RECT  52.12 110.85 52.77 110.99 ;
      RECT  52.96 110.86 53.68 111.0 ;
      RECT  52.12 110.99 52.26 115.88 ;
      RECT  53.54 110.14 53.68 110.86 ;
      RECT  53.54 111.0 53.68 115.88 ;
      RECT  52.45 120.33 52.77 120.22 ;
      RECT  52.96 120.32 53.28 120.22 ;
      RECT  52.45 120.54 52.77 120.47 ;
      RECT  52.96 120.54 53.28 120.46 ;
      RECT  52.12 121.18 52.26 120.47 ;
      RECT  52.12 120.47 52.77 120.33 ;
      RECT  52.96 120.46 53.68 120.32 ;
      RECT  52.12 120.33 52.26 115.44 ;
      RECT  53.54 121.18 53.68 120.46 ;
      RECT  53.54 120.32 53.68 115.44 ;
      RECT  52.12 120.78 52.26 126.52 ;
      RECT  53.54 120.78 53.68 126.52 ;
      RECT  52.12 25.22 52.26 126.3 ;
      RECT  53.54 25.22 53.68 126.3 ;
      RECT  56.12 36.06 56.26 30.32 ;
      RECT  57.54 36.06 57.68 30.32 ;
      RECT  60.12 36.06 60.26 30.32 ;
      RECT  61.54 36.06 61.68 30.32 ;
      RECT  56.12 35.86 56.26 30.54 ;
      RECT  57.54 35.86 57.68 30.54 ;
      RECT  60.12 35.86 60.26 30.54 ;
      RECT  61.54 35.86 61.68 30.54 ;
      RECT  56.12 25.02 56.26 30.76 ;
      RECT  57.54 25.02 57.68 30.76 ;
      RECT  60.12 25.02 60.26 30.76 ;
      RECT  61.54 25.02 61.68 30.76 ;
      RECT  56.12 25.22 56.26 30.54 ;
      RECT  57.54 25.22 57.68 30.54 ;
      RECT  60.12 25.22 60.26 30.54 ;
      RECT  61.54 25.22 61.68 30.54 ;
      RECT  56.12 120.78 56.26 126.52 ;
      RECT  57.54 120.78 57.68 126.52 ;
      RECT  60.12 120.78 60.26 126.52 ;
      RECT  61.54 120.78 61.68 126.52 ;
      RECT  56.12 120.98 56.26 126.3 ;
      RECT  57.54 120.98 57.68 126.3 ;
      RECT  60.12 120.98 60.26 126.3 ;
      RECT  61.54 120.98 61.68 126.3 ;
      RECT  48.12 25.02 48.26 30.76 ;
      RECT  49.54 25.02 49.68 30.76 ;
      RECT  48.12 36.06 48.26 30.32 ;
      RECT  49.54 36.06 49.68 30.32 ;
      RECT  48.12 35.66 48.26 41.4 ;
      RECT  49.54 35.66 49.68 41.4 ;
      RECT  48.12 46.7 48.26 40.96 ;
      RECT  49.54 46.7 49.68 40.96 ;
      RECT  48.12 46.3 48.26 52.04 ;
      RECT  49.54 46.3 49.68 52.04 ;
      RECT  48.12 57.34 48.26 51.6 ;
      RECT  49.54 57.34 49.68 51.6 ;
      RECT  48.12 56.94 48.26 62.68 ;
      RECT  49.54 56.94 49.68 62.68 ;
      RECT  48.12 67.98 48.26 62.24 ;
      RECT  49.54 67.98 49.68 62.24 ;
      RECT  48.12 67.58 48.26 73.32 ;
      RECT  49.54 67.58 49.68 73.32 ;
      RECT  48.12 78.62 48.26 72.88 ;
      RECT  49.54 78.62 49.68 72.88 ;
      RECT  48.12 78.22 48.26 83.96 ;
      RECT  49.54 78.22 49.68 83.96 ;
      RECT  48.12 89.26 48.26 83.52 ;
      RECT  49.54 89.26 49.68 83.52 ;
      RECT  48.12 88.86 48.26 94.6 ;
      RECT  49.54 88.86 49.68 94.6 ;
      RECT  48.12 99.9 48.26 94.16 ;
      RECT  49.54 99.9 49.68 94.16 ;
      RECT  48.12 99.5 48.26 105.24 ;
      RECT  49.54 99.5 49.68 105.24 ;
      RECT  48.12 110.54 48.26 104.8 ;
      RECT  49.54 110.54 49.68 104.8 ;
      RECT  48.12 110.14 48.26 115.88 ;
      RECT  49.54 110.14 49.68 115.88 ;
      RECT  48.12 121.18 48.26 115.44 ;
      RECT  49.54 121.18 49.68 115.44 ;
      RECT  48.12 120.78 48.26 126.52 ;
      RECT  49.54 120.78 49.68 126.52 ;
      RECT  48.12 25.22 48.26 126.3 ;
      RECT  49.54 25.22 49.68 126.3 ;
      RECT  64.12 25.02 64.26 30.76 ;
      RECT  65.54 25.02 65.68 30.76 ;
      RECT  64.12 36.06 64.26 30.32 ;
      RECT  65.54 36.06 65.68 30.32 ;
      RECT  64.12 35.66 64.26 41.4 ;
      RECT  65.54 35.66 65.68 41.4 ;
      RECT  64.12 46.7 64.26 40.96 ;
      RECT  65.54 46.7 65.68 40.96 ;
      RECT  64.12 46.3 64.26 52.04 ;
      RECT  65.54 46.3 65.68 52.04 ;
      RECT  64.12 57.34 64.26 51.6 ;
      RECT  65.54 57.34 65.68 51.6 ;
      RECT  64.12 56.94 64.26 62.68 ;
      RECT  65.54 56.94 65.68 62.68 ;
      RECT  64.12 67.98 64.26 62.24 ;
      RECT  65.54 67.98 65.68 62.24 ;
      RECT  64.12 67.58 64.26 73.32 ;
      RECT  65.54 67.58 65.68 73.32 ;
      RECT  64.12 78.62 64.26 72.88 ;
      RECT  65.54 78.62 65.68 72.88 ;
      RECT  64.12 78.22 64.26 83.96 ;
      RECT  65.54 78.22 65.68 83.96 ;
      RECT  64.12 89.26 64.26 83.52 ;
      RECT  65.54 89.26 65.68 83.52 ;
      RECT  64.12 88.86 64.26 94.6 ;
      RECT  65.54 88.86 65.68 94.6 ;
      RECT  64.12 99.9 64.26 94.16 ;
      RECT  65.54 99.9 65.68 94.16 ;
      RECT  64.12 99.5 64.26 105.24 ;
      RECT  65.54 99.5 65.68 105.24 ;
      RECT  64.12 110.54 64.26 104.8 ;
      RECT  65.54 110.54 65.68 104.8 ;
      RECT  64.12 110.14 64.26 115.88 ;
      RECT  65.54 110.14 65.68 115.88 ;
      RECT  64.12 121.18 64.26 115.44 ;
      RECT  65.54 121.18 65.68 115.44 ;
      RECT  64.12 120.78 64.26 126.52 ;
      RECT  65.54 120.78 65.68 126.52 ;
      RECT  64.12 25.22 64.26 126.3 ;
      RECT  65.54 25.22 65.68 126.3 ;
      RECT  52.12 25.22 52.26 126.3 ;
      RECT  53.54 25.22 53.68 126.3 ;
      RECT  56.12 25.22 56.77 126.3 ;
      RECT  56.96 25.22 57.68 126.3 ;
      RECT  60.12 25.22 60.77 126.3 ;
      RECT  60.96 25.22 61.68 126.3 ;
      RECT  51.52 15.82 51.66 23.12 ;
      RECT  54.12 15.82 54.26 23.12 ;
      RECT  55.52 15.82 55.66 23.12 ;
      RECT  58.12 15.82 58.26 23.12 ;
      RECT  59.52 15.82 59.66 23.12 ;
      RECT  62.12 15.82 62.26 23.12 ;
      RECT  51.52 15.82 51.66 23.12 ;
      RECT  54.12 15.82 54.26 23.12 ;
      RECT  55.52 15.82 55.66 23.12 ;
      RECT  58.12 15.82 58.26 23.12 ;
      RECT  59.52 15.82 59.66 23.12 ;
      RECT  62.12 15.82 62.26 23.12 ;
      RECT  56.39 11.23 56.72 11.56 ;
      RECT  56.39 11.56 56.53 14.17 ;
      RECT  57.5 9.06 57.64 10.61 ;
      RECT  56.39 9.06 56.53 11.23 ;
      RECT  58.05 13.5 58.5 13.95 ;
      RECT  58.19 9.04 58.64 9.49 ;
      RECT  57.5 10.61 57.96 10.94 ;
      RECT  57.5 10.94 57.64 14.17 ;
      RECT  60.39 11.23 60.72 11.56 ;
      RECT  60.39 11.56 60.53 14.17 ;
      RECT  61.5 9.06 61.64 10.61 ;
      RECT  60.39 9.06 60.53 11.23 ;
      RECT  62.05 13.5 62.5 13.95 ;
      RECT  62.19 9.04 62.64 9.49 ;
      RECT  61.5 10.61 61.96 10.94 ;
      RECT  61.5 10.94 61.64 14.17 ;
      RECT  56.39 11.23 56.72 11.56 ;
      RECT  57.5 10.61 57.96 10.94 ;
      RECT  60.39 11.23 60.72 11.56 ;
      RECT  61.5 10.61 61.96 10.94 ;
      RECT  51.52 23.12 51.66 15.82 ;
      RECT  54.12 23.12 54.26 15.82 ;
      RECT  55.52 23.12 55.66 15.82 ;
      RECT  58.12 23.12 58.26 15.82 ;
      RECT  59.52 23.12 59.66 15.82 ;
      RECT  62.12 23.12 62.26 15.82 ;
      RECT  3.74 38.18 4.2 38.64 ;
      RECT  4.44 43.72 4.9 44.18 ;
      RECT  3.74 70.1 4.2 70.56 ;
      RECT  4.44 75.64 4.9 76.1 ;
      RECT  0.16 35.86 0.3 89.06 ;
      RECT  0.86 35.86 1.0 89.06 ;
      RECT  1.56 35.86 1.7 89.06 ;
      RECT  2.26 35.86 2.4 89.06 ;
      RECT  37.41 35.86 37.55 120.98 ;
      RECT  0.16 35.86 0.3 89.06 ;
      RECT  0.86 35.86 1.0 89.06 ;
      RECT  1.56 35.86 1.7 89.06 ;
      RECT  2.26 35.86 2.4 89.06 ;
      RECT  36.82 34.37 36.96 34.51 ;
      RECT  0.16 35.86 0.3 89.06 ;
      RECT  0.86 35.86 1.0 89.06 ;
      RECT  1.56 35.86 1.7 89.06 ;
      RECT  2.26 35.86 2.4 89.06 ;
      RECT  40.53 0.0 40.67 25.22 ;
      RECT  42.35 0.0 42.49 25.22 ;
      RECT  41.44 0.0 41.58 25.22 ;
      RECT  43.26 0.0 43.4 25.22 ;
      RECT  -52.59 -8.52 -52.28 -8.2 ;
      RECT  -42.54 -7.96 -42.22 -7.64 ;
      RECT  -51.1 -7.28 -50.76 -6.96 ;
      RECT  -51.1 -7.28 -50.76 -6.96 ;
      RECT  -29.76 -9.54 -29.62 -9.4 ;
      RECT  -33.35 -6.71 -33.21 -6.57 ;
      RECT  -52.59 -8.52 -52.28 -8.2 ;
      RECT  -52.59 -3.08 -52.28 -3.4 ;
      RECT  -42.54 -3.64 -42.22 -3.96 ;
      RECT  -51.1 -4.32 -50.76 -4.64 ;
      RECT  -51.1 -4.32 -50.76 -4.64 ;
      RECT  -29.76 -2.06 -29.62 -2.2 ;
      RECT  -33.35 -4.89 -33.21 -5.03 ;
      RECT  -52.59 -3.08 -52.28 -3.4 ;
      RECT  -51.1 -7.28 -50.76 -6.96 ;
      RECT  -51.1 -4.64 -50.76 -4.32 ;
      RECT  -29.76 -9.54 -29.62 -9.4 ;
      RECT  -33.35 -6.71 -33.21 -6.57 ;
      RECT  -29.76 -2.2 -29.62 -2.06 ;
      RECT  -33.35 -5.03 -33.21 -4.89 ;
      RECT  -52.59 -10.06 -52.45 -1.54 ;
      RECT  -37.1 25.22 -37.24 29.31 ;
      RECT  -51.33 25.22 -51.47 96.51 ;
      RECT  -51.1 -7.28 -50.76 -6.96 ;
      RECT  -51.1 -4.64 -50.76 -4.32 ;
      RECT  -20.88 -8.11 -20.74 -7.97 ;
      RECT  -37.24 25.22 -37.1 29.31 ;
      RECT  -15.16 21.93 -1.4 22.07 ;
      RECT  -14.08 8.87 -1.4 9.01 ;
      RECT  -12.54 13.41 -1.4 13.55 ;
      RECT  -8.34 4.95 -1.4 5.09 ;
      RECT  -5.64 -8.17 -1.4 -8.03 ;
      RECT  -14.28 103.56 -13.97 103.88 ;
      RECT  -4.23 104.12 -3.91 104.44 ;
      RECT  -12.79 104.8 -12.45 105.12 ;
      RECT  -14.28 109.0 -13.97 108.68 ;
      RECT  -4.23 108.44 -3.91 108.12 ;
      RECT  -12.79 107.76 -12.45 107.44 ;
      RECT  -14.28 112.08 -13.97 112.4 ;
      RECT  -4.23 112.64 -3.91 112.96 ;
      RECT  -12.79 113.32 -12.45 113.64 ;
      RECT  -14.28 117.52 -13.97 117.2 ;
      RECT  -4.23 116.96 -3.91 116.64 ;
      RECT  -12.79 116.28 -12.45 115.96 ;
      RECT  -12.79 104.8 -12.45 105.12 ;
      RECT  -12.79 107.44 -12.45 107.76 ;
      RECT  -12.79 113.32 -12.45 113.64 ;
      RECT  -12.79 115.96 -12.45 116.28 ;
      RECT  -4.23 104.12 -3.91 104.44 ;
      RECT  -4.23 108.12 -3.91 108.44 ;
      RECT  -4.23 112.64 -3.91 112.96 ;
      RECT  -4.23 116.64 -3.91 116.96 ;
      RECT  11.98 -8.52 12.29 -8.2 ;
      RECT  22.03 -7.96 22.35 -7.64 ;
      RECT  13.47 -7.28 13.81 -6.96 ;
      RECT  25.11 -8.52 25.42 -8.2 ;
      RECT  35.16 -7.96 35.48 -7.64 ;
      RECT  26.6 -7.28 26.94 -6.96 ;
      RECT  13.47 -7.28 13.81 -6.96 ;
      RECT  26.6 -7.28 26.94 -6.96 ;
      RECT  22.03 -7.96 22.35 -7.64 ;
      RECT  35.16 -7.96 35.48 -7.64 ;
   LAYER  m3 ;
      RECT  52.66 30.3 53.12 30.76 ;
      RECT  52.66 126.06 53.12 126.52 ;
      RECT  52.66 120.76 53.12 121.22 ;
      RECT  52.66 25.0 53.12 25.46 ;
      RECT  48.66 104.8 49.12 105.26 ;
      RECT  64.66 83.5 65.12 83.96 ;
      RECT  64.66 40.96 65.12 41.42 ;
      RECT  64.66 62.24 65.12 62.7 ;
      RECT  64.66 62.22 65.12 62.68 ;
      RECT  64.66 51.58 65.12 52.04 ;
      RECT  52.66 126.06 53.12 126.52 ;
      RECT  48.66 72.86 49.12 73.32 ;
      RECT  64.66 30.32 65.12 30.78 ;
      RECT  64.66 104.78 65.12 105.24 ;
      RECT  64.66 72.86 65.12 73.32 ;
      RECT  48.66 40.96 49.12 41.42 ;
      RECT  48.66 62.24 49.12 62.7 ;
      RECT  64.66 94.14 65.12 94.6 ;
      RECT  52.66 30.3 53.12 30.76 ;
      RECT  48.66 104.78 49.12 105.24 ;
      RECT  64.66 94.16 65.12 94.62 ;
      RECT  48.66 83.52 49.12 83.98 ;
      RECT  48.66 40.94 49.12 41.4 ;
      RECT  48.66 83.5 49.12 83.96 ;
      RECT  64.66 51.6 65.12 52.06 ;
      RECT  48.66 30.3 49.12 30.76 ;
      RECT  48.66 94.16 49.12 94.62 ;
      RECT  60.66 126.06 61.12 126.52 ;
      RECT  64.66 126.06 65.12 126.52 ;
      RECT  48.66 62.22 49.12 62.68 ;
      RECT  64.66 40.94 65.12 41.4 ;
      RECT  48.66 115.42 49.12 115.88 ;
      RECT  56.66 30.3 57.12 30.76 ;
      RECT  48.66 94.14 49.12 94.6 ;
      RECT  64.66 115.44 65.12 115.9 ;
      RECT  56.66 126.06 57.12 126.52 ;
      RECT  64.66 115.42 65.12 115.88 ;
      RECT  60.66 30.3 61.12 30.76 ;
      RECT  48.66 51.6 49.12 52.06 ;
      RECT  48.66 30.32 49.12 30.78 ;
      RECT  48.66 51.58 49.12 52.04 ;
      RECT  64.66 30.3 65.12 30.76 ;
      RECT  48.66 126.06 49.12 126.52 ;
      RECT  48.66 72.88 49.12 73.34 ;
      RECT  64.66 83.52 65.12 83.98 ;
      RECT  64.66 104.8 65.12 105.26 ;
      RECT  48.66 115.44 49.12 115.9 ;
      RECT  64.66 72.88 65.12 73.34 ;
      RECT  48.66 56.9 49.12 57.36 ;
      RECT  48.66 46.28 49.12 46.74 ;
      RECT  64.66 110.1 65.12 110.56 ;
      RECT  64.66 99.46 65.12 99.92 ;
      RECT  64.66 110.12 65.12 110.58 ;
      RECT  60.66 120.76 61.12 121.22 ;
      RECT  64.66 46.28 65.12 46.74 ;
      RECT  64.66 120.76 65.12 121.22 ;
      RECT  52.66 120.76 53.12 121.22 ;
      RECT  64.66 67.54 65.12 68.0 ;
      RECT  67.56 26.14 68.02 26.6 ;
      RECT  67.56 121.9 68.02 122.36 ;
      RECT  48.66 88.82 49.12 89.28 ;
      RECT  48.66 120.76 49.12 121.22 ;
      RECT  48.66 120.74 49.12 121.2 ;
      RECT  48.66 99.46 49.12 99.92 ;
      RECT  48.66 56.92 49.12 57.38 ;
      RECT  64.66 67.56 65.12 68.02 ;
      RECT  60.66 25.0 61.12 25.46 ;
      RECT  48.66 35.62 49.12 36.08 ;
      RECT  64.66 88.82 65.12 89.28 ;
      RECT  64.66 99.48 65.12 99.94 ;
      RECT  48.66 110.12 49.12 110.58 ;
      RECT  48.66 78.2 49.12 78.66 ;
      RECT  48.66 67.54 49.12 68.0 ;
      RECT  64.66 46.26 65.12 46.72 ;
      RECT  64.66 56.9 65.12 57.36 ;
      RECT  56.66 120.76 57.12 121.22 ;
      RECT  64.66 25.0 65.12 25.46 ;
      RECT  48.66 67.56 49.12 68.02 ;
      RECT  52.66 25.0 53.12 25.46 ;
      RECT  64.66 35.64 65.12 36.1 ;
      RECT  64.66 88.84 65.12 89.3 ;
      RECT  45.76 26.14 46.22 26.6 ;
      RECT  45.76 121.9 46.22 122.36 ;
      RECT  48.66 78.18 49.12 78.64 ;
      RECT  64.66 56.92 65.12 57.38 ;
      RECT  64.66 120.74 65.12 121.2 ;
      RECT  64.66 78.2 65.12 78.66 ;
      RECT  48.66 110.1 49.12 110.56 ;
      RECT  64.66 35.62 65.12 36.08 ;
      RECT  48.66 99.48 49.12 99.94 ;
      RECT  56.66 25.0 57.12 25.46 ;
      RECT  48.66 25.0 49.12 25.46 ;
      RECT  48.66 35.64 49.12 36.1 ;
      RECT  64.66 78.18 65.12 78.64 ;
      RECT  48.66 88.84 49.12 89.3 ;
      RECT  48.66 46.26 49.12 46.72 ;
      RECT  52.89 22.33 53.35 22.79 ;
      RECT  56.89 22.33 57.35 22.79 ;
      RECT  60.89 22.33 61.35 22.79 ;
      RECT  60.89 22.33 61.35 22.79 ;
      RECT  56.89 22.33 57.35 22.79 ;
      RECT  52.89 22.33 53.35 22.79 ;
      RECT  57.99 13.47 58.52 13.97 ;
      RECT  58.14 9.02 58.66 9.52 ;
      RECT  61.99 13.47 62.52 13.97 ;
      RECT  62.14 9.02 62.66 9.52 ;
      RECT  56.66 13.49 57.12 13.95 ;
      RECT  60.66 13.49 61.12 13.95 ;
      RECT  60.66 9.03 61.12 9.49 ;
      RECT  56.66 9.03 57.12 9.49 ;
      RECT  65.95 6.94 66.41 7.4 ;
      RECT  61.95 6.94 62.41 7.4 ;
      RECT  61.95 1.13 62.41 1.59 ;
      RECT  65.95 1.13 66.41 1.59 ;
      RECT  56.89 22.79 57.35 22.33 ;
      RECT  52.89 22.79 53.35 22.33 ;
      RECT  60.89 22.79 61.35 22.33 ;
      RECT  56.66 13.95 57.12 13.49 ;
      RECT  61.95 7.4 62.41 6.94 ;
      RECT  60.66 13.95 61.12 13.49 ;
      RECT  65.95 7.4 66.41 6.94 ;
      RECT  56.66 9.49 57.12 9.03 ;
      RECT  61.95 1.59 62.41 1.13 ;
      RECT  60.66 9.49 61.12 9.03 ;
      RECT  65.95 1.59 66.41 1.13 ;
      RECT  5.53 51.59 5.99 52.05 ;
      RECT  13.16 51.59 13.62 52.05 ;
      RECT  5.53 40.95 5.99 41.41 ;
      RECT  13.16 40.95 13.62 41.41 ;
      RECT  5.53 56.91 5.99 57.37 ;
      RECT  5.53 35.63 5.99 36.09 ;
      RECT  13.16 35.63 13.62 36.09 ;
      RECT  13.16 56.91 13.62 57.37 ;
      RECT  13.16 46.27 13.62 46.73 ;
      RECT  5.53 46.27 5.99 46.73 ;
      RECT  5.53 83.51 5.99 83.97 ;
      RECT  13.16 83.51 13.62 83.97 ;
      RECT  5.53 72.87 5.99 73.33 ;
      RECT  13.16 72.87 13.62 73.33 ;
      RECT  5.53 88.83 5.99 89.29 ;
      RECT  5.53 67.55 5.99 68.01 ;
      RECT  13.16 67.55 13.62 68.01 ;
      RECT  13.16 88.83 13.62 89.29 ;
      RECT  13.16 78.19 13.62 78.65 ;
      RECT  5.53 78.19 5.99 78.65 ;
      RECT  34.85 72.87 35.31 73.33 ;
      RECT  34.85 104.79 35.31 105.25 ;
      RECT  34.85 104.79 35.31 105.25 ;
      RECT  34.85 94.15 35.31 94.61 ;
      RECT  5.53 51.59 5.99 52.05 ;
      RECT  34.85 40.95 35.31 41.41 ;
      RECT  34.85 83.51 35.31 83.97 ;
      RECT  34.85 51.59 35.31 52.05 ;
      RECT  34.85 115.43 35.31 115.89 ;
      RECT  34.85 115.43 35.31 115.89 ;
      RECT  13.16 51.59 13.62 52.05 ;
      RECT  5.53 40.95 5.99 41.41 ;
      RECT  5.53 83.51 5.99 83.97 ;
      RECT  13.16 83.51 13.62 83.97 ;
      RECT  13.16 40.95 13.62 41.41 ;
      RECT  13.16 72.87 13.62 73.33 ;
      RECT  34.85 62.23 35.31 62.69 ;
      RECT  5.53 72.87 5.99 73.33 ;
      RECT  5.53 56.91 5.99 57.37 ;
      RECT  5.53 88.83 5.99 89.29 ;
      RECT  13.16 56.91 13.62 57.37 ;
      RECT  5.53 67.55 5.99 68.01 ;
      RECT  5.53 46.27 5.99 46.73 ;
      RECT  13.16 88.83 13.62 89.29 ;
      RECT  13.16 78.19 13.62 78.65 ;
      RECT  34.85 120.75 35.31 121.21 ;
      RECT  34.85 110.11 35.31 110.57 ;
      RECT  34.85 46.27 35.31 46.73 ;
      RECT  34.85 78.19 35.31 78.65 ;
      RECT  13.16 46.27 13.62 46.73 ;
      RECT  34.85 88.83 35.31 89.29 ;
      RECT  5.53 78.19 5.99 78.65 ;
      RECT  34.85 99.47 35.31 99.93 ;
      RECT  34.85 67.55 35.31 68.01 ;
      RECT  5.53 35.63 5.99 36.09 ;
      RECT  13.16 35.63 13.62 36.09 ;
      RECT  34.85 35.63 35.31 36.09 ;
      RECT  13.16 67.55 13.62 68.01 ;
      RECT  34.85 56.91 35.31 57.37 ;
      RECT  42.39 51.59 42.85 52.05 ;
      RECT  42.39 104.79 42.85 105.25 ;
      RECT  42.39 104.79 42.85 105.25 ;
      RECT  42.39 115.43 42.85 115.89 ;
      RECT  42.39 115.43 42.85 115.89 ;
      RECT  42.39 94.15 42.85 94.61 ;
      RECT  42.39 83.51 42.85 83.97 ;
      RECT  42.39 62.23 42.85 62.69 ;
      RECT  42.39 40.95 42.85 41.41 ;
      RECT  42.39 72.87 42.85 73.33 ;
      RECT  42.39 78.19 42.85 78.65 ;
      RECT  42.39 99.47 42.85 99.93 ;
      RECT  42.39 110.11 42.85 110.57 ;
      RECT  42.39 120.75 42.85 121.21 ;
      RECT  42.39 35.63 42.85 36.09 ;
      RECT  42.39 67.55 42.85 68.01 ;
      RECT  42.39 56.91 42.85 57.37 ;
      RECT  42.39 88.83 42.85 89.29 ;
      RECT  42.39 46.27 42.85 46.73 ;
      RECT  42.39 40.95 42.85 41.41 ;
      RECT  42.39 51.59 42.85 52.05 ;
      RECT  42.39 62.23 42.85 62.69 ;
      RECT  42.39 104.79 42.85 105.25 ;
      RECT  35.54 32.39 36.0 32.85 ;
      RECT  5.53 72.87 5.99 73.33 ;
      RECT  34.85 115.43 35.31 115.89 ;
      RECT  5.53 83.51 5.99 83.97 ;
      RECT  34.85 51.59 35.31 52.05 ;
      RECT  5.53 40.95 5.99 41.41 ;
      RECT  13.16 83.51 13.62 83.97 ;
      RECT  34.85 72.87 35.31 73.33 ;
      RECT  13.16 51.59 13.62 52.05 ;
      RECT  42.39 83.51 42.85 83.97 ;
      RECT  34.85 104.79 35.31 105.25 ;
      RECT  34.85 62.23 35.31 62.69 ;
      RECT  42.39 115.43 42.85 115.89 ;
      RECT  34.85 94.15 35.31 94.61 ;
      RECT  13.16 40.95 13.62 41.41 ;
      RECT  34.85 30.31 35.31 30.77 ;
      RECT  34.85 40.95 35.31 41.41 ;
      RECT  42.39 94.15 42.85 94.61 ;
      RECT  13.16 72.87 13.62 73.33 ;
      RECT  42.39 72.87 42.85 73.33 ;
      RECT  5.53 51.59 5.99 52.05 ;
      RECT  34.85 83.51 35.31 83.97 ;
      RECT  42.39 56.91 42.85 57.37 ;
      RECT  13.16 67.55 13.62 68.01 ;
      RECT  5.53 88.83 5.99 89.29 ;
      RECT  5.53 35.63 5.99 36.09 ;
      RECT  34.85 35.63 35.31 36.09 ;
      RECT  13.16 35.63 13.62 36.09 ;
      RECT  5.53 56.91 5.99 57.37 ;
      RECT  34.85 78.19 35.31 78.65 ;
      RECT  13.16 46.27 13.62 46.73 ;
      RECT  13.16 56.91 13.62 57.37 ;
      RECT  42.39 78.19 42.85 78.65 ;
      RECT  42.39 46.27 42.85 46.73 ;
      RECT  34.85 120.75 35.31 121.21 ;
      RECT  34.85 67.55 35.31 68.01 ;
      RECT  42.39 120.75 42.85 121.21 ;
      RECT  42.39 99.47 42.85 99.93 ;
      RECT  5.53 67.55 5.99 68.01 ;
      RECT  42.39 88.83 42.85 89.29 ;
      RECT  42.39 35.63 42.85 36.09 ;
      RECT  13.16 78.19 13.62 78.65 ;
      RECT  13.16 88.83 13.62 89.29 ;
      RECT  34.85 99.47 35.31 99.93 ;
      RECT  42.39 110.11 42.85 110.57 ;
      RECT  5.53 46.27 5.99 46.73 ;
      RECT  34.85 110.11 35.31 110.57 ;
      RECT  34.85 46.27 35.31 46.73 ;
      RECT  34.85 88.83 35.31 89.29 ;
      RECT  5.53 78.19 5.99 78.65 ;
      RECT  42.39 67.55 42.85 68.01 ;
      RECT  34.85 56.91 35.31 57.37 ;
      RECT  0.0 14.76 51.59 15.06 ;
      RECT  64.66 83.5 65.12 83.96 ;
      RECT  34.85 115.43 35.31 115.89 ;
      RECT  64.66 104.78 65.12 105.24 ;
      RECT  48.66 62.24 49.12 62.7 ;
      RECT  64.66 51.6 65.12 52.06 ;
      RECT  42.39 104.79 42.85 105.25 ;
      RECT  56.89 22.33 57.35 22.79 ;
      RECT  48.66 62.22 49.12 62.68 ;
      RECT  64.66 115.44 65.12 115.9 ;
      RECT  60.66 30.3 61.12 30.76 ;
      RECT  48.66 126.06 49.12 126.52 ;
      RECT  64.66 83.52 65.12 83.98 ;
      RECT  42.39 40.95 42.85 41.41 ;
      RECT  64.66 40.96 65.12 41.42 ;
      RECT  52.66 126.06 53.12 126.52 ;
      RECT  64.66 30.32 65.12 30.78 ;
      RECT  13.16 40.95 13.62 41.41 ;
      RECT  34.85 94.15 35.31 94.61 ;
      RECT  5.53 83.51 5.99 83.97 ;
      RECT  48.66 104.78 49.12 105.24 ;
      RECT  48.66 40.94 49.12 41.4 ;
      RECT  48.66 83.5 49.12 83.96 ;
      RECT  34.85 51.59 35.31 52.05 ;
      RECT  48.66 94.16 49.12 94.62 ;
      RECT  60.66 126.06 61.12 126.52 ;
      RECT  34.85 83.51 35.31 83.97 ;
      RECT  48.66 94.14 49.12 94.6 ;
      RECT  56.66 126.06 57.12 126.52 ;
      RECT  48.66 51.6 49.12 52.06 ;
      RECT  52.89 22.33 53.35 22.79 ;
      RECT  64.66 30.3 65.12 30.76 ;
      RECT  13.16 72.87 13.62 73.33 ;
      RECT  48.66 115.44 49.12 115.9 ;
      RECT  64.66 72.88 65.12 73.34 ;
      RECT  61.95 6.94 62.41 7.4 ;
      RECT  64.66 62.24 65.12 62.7 ;
      RECT  64.66 51.58 65.12 52.04 ;
      RECT  48.66 72.86 49.12 73.32 ;
      RECT  64.66 72.86 65.12 73.32 ;
      RECT  48.66 40.96 49.12 41.42 ;
      RECT  35.54 32.39 36.0 32.85 ;
      RECT  64.66 94.16 65.12 94.62 ;
      RECT  42.39 83.51 42.85 83.97 ;
      RECT  56.66 13.49 57.12 13.95 ;
      RECT  60.89 22.33 61.35 22.79 ;
      RECT  5.53 72.87 5.99 73.33 ;
      RECT  64.66 40.94 65.12 41.4 ;
      RECT  5.53 51.59 5.99 52.05 ;
      RECT  48.66 115.42 49.12 115.88 ;
      RECT  34.85 62.23 35.31 62.69 ;
      RECT  64.66 115.42 65.12 115.88 ;
      RECT  34.85 104.79 35.31 105.25 ;
      RECT  48.66 51.58 49.12 52.04 ;
      RECT  42.39 51.59 42.85 52.05 ;
      RECT  13.16 83.51 13.62 83.97 ;
      RECT  48.66 104.8 49.12 105.26 ;
      RECT  13.16 51.59 13.62 52.05 ;
      RECT  42.39 72.87 42.85 73.33 ;
      RECT  5.53 40.95 5.99 41.41 ;
      RECT  42.39 62.23 42.85 62.69 ;
      RECT  64.66 62.22 65.12 62.68 ;
      RECT  34.85 30.31 35.31 30.77 ;
      RECT  64.66 94.14 65.12 94.6 ;
      RECT  34.85 72.87 35.31 73.33 ;
      RECT  52.66 30.3 53.12 30.76 ;
      RECT  48.66 83.52 49.12 83.98 ;
      RECT  48.66 30.3 49.12 30.76 ;
      RECT  42.39 94.15 42.85 94.61 ;
      RECT  64.66 126.06 65.12 126.52 ;
      RECT  34.85 40.95 35.31 41.41 ;
      RECT  56.66 30.3 57.12 30.76 ;
      RECT  60.66 13.49 61.12 13.95 ;
      RECT  48.66 30.32 49.12 30.78 ;
      RECT  48.66 72.88 49.12 73.34 ;
      RECT  64.66 104.8 65.12 105.26 ;
      RECT  65.95 6.94 66.41 7.4 ;
      RECT  42.39 115.43 42.85 115.89 ;
      RECT  48.66 56.9 49.12 57.36 ;
      RECT  48.66 46.28 49.12 46.74 ;
      RECT  34.85 35.63 35.31 36.09 ;
      RECT  34.85 46.27 35.31 46.73 ;
      RECT  64.66 46.28 65.12 46.74 ;
      RECT  42.39 35.63 42.85 36.09 ;
      RECT  34.85 88.83 35.31 89.29 ;
      RECT  60.66 9.03 61.12 9.49 ;
      RECT  64.66 67.54 65.12 68.0 ;
      RECT  48.66 120.74 49.12 121.2 ;
      RECT  48.66 99.46 49.12 99.92 ;
      RECT  60.66 25.0 61.12 25.46 ;
      RECT  48.66 35.62 49.12 36.08 ;
      RECT  64.66 35.64 65.12 36.1 ;
      RECT  64.66 56.92 65.12 57.38 ;
      RECT  64.66 120.74 65.12 121.2 ;
      RECT  64.66 78.2 65.12 78.66 ;
      RECT  48.66 110.1 49.12 110.56 ;
      RECT  48.66 99.48 49.12 99.94 ;
      RECT  56.66 25.0 57.12 25.46 ;
      RECT  48.66 35.64 49.12 36.1 ;
      RECT  48.66 88.84 49.12 89.3 ;
      RECT  56.66 9.03 57.12 9.49 ;
      RECT  64.66 110.1 65.12 110.56 ;
      RECT  64.66 110.12 65.12 110.58 ;
      RECT  67.56 121.9 68.02 122.36 ;
      RECT  5.53 88.83 5.99 89.29 ;
      RECT  48.66 88.82 49.12 89.28 ;
      RECT  5.53 56.91 5.99 57.37 ;
      RECT  13.16 46.27 13.62 46.73 ;
      RECT  34.85 78.19 35.31 78.65 ;
      RECT  34.85 67.55 35.31 68.01 ;
      RECT  34.85 56.91 35.31 57.37 ;
      RECT  48.66 78.2 49.12 78.66 ;
      RECT  64.66 46.26 65.12 46.72 ;
      RECT  48.66 67.54 49.12 68.0 ;
      RECT  56.66 120.76 57.12 121.22 ;
      RECT  65.95 1.13 66.41 1.59 ;
      RECT  42.39 78.19 42.85 78.65 ;
      RECT  45.76 121.9 46.22 122.36 ;
      RECT  48.66 78.18 49.12 78.64 ;
      RECT  48.66 46.26 49.12 46.72 ;
      RECT  34.85 99.47 35.31 99.93 ;
      RECT  13.16 67.55 13.62 68.01 ;
      RECT  64.66 99.46 65.12 99.92 ;
      RECT  60.66 120.76 61.12 121.22 ;
      RECT  52.66 120.76 53.12 121.22 ;
      RECT  67.56 26.14 68.02 26.6 ;
      RECT  48.66 120.76 49.12 121.22 ;
      RECT  34.85 120.75 35.31 121.21 ;
      RECT  5.53 78.19 5.99 78.65 ;
      RECT  61.95 1.13 62.41 1.59 ;
      RECT  64.66 88.82 65.12 89.28 ;
      RECT  64.66 99.48 65.12 99.94 ;
      RECT  48.66 110.12 49.12 110.58 ;
      RECT  64.66 25.0 65.12 25.46 ;
      RECT  48.66 67.56 49.12 68.02 ;
      RECT  5.53 35.63 5.99 36.09 ;
      RECT  42.39 56.91 42.85 57.37 ;
      RECT  13.16 35.63 13.62 36.09 ;
      RECT  42.39 67.55 42.85 68.01 ;
      RECT  13.16 56.91 13.62 57.37 ;
      RECT  48.66 25.0 49.12 25.46 ;
      RECT  64.66 78.18 65.12 78.64 ;
      RECT  42.39 88.83 42.85 89.29 ;
      RECT  42.39 120.75 42.85 121.21 ;
      RECT  42.39 46.27 42.85 46.73 ;
      RECT  13.16 78.19 13.62 78.65 ;
      RECT  64.66 120.76 65.12 121.22 ;
      RECT  5.53 46.27 5.99 46.73 ;
      RECT  48.66 56.92 49.12 57.38 ;
      RECT  64.66 67.56 65.12 68.02 ;
      RECT  34.85 110.11 35.31 110.57 ;
      RECT  5.53 67.55 5.99 68.01 ;
      RECT  64.66 56.9 65.12 57.36 ;
      RECT  52.66 25.0 53.12 25.46 ;
      RECT  64.66 88.84 65.12 89.3 ;
      RECT  45.76 26.14 46.22 26.6 ;
      RECT  42.39 99.47 42.85 99.93 ;
      RECT  13.16 88.83 13.62 89.29 ;
      RECT  64.66 35.62 65.12 36.08 ;
      RECT  42.39 110.11 42.85 110.57 ;
      RECT  -53.07 -6.02 -52.61 -5.56 ;
      RECT  -53.07 -6.04 -52.61 -5.58 ;
      RECT  -53.07 -1.8 -52.61 -1.34 ;
      RECT  -53.07 -10.26 -52.61 -9.8 ;
      RECT  -48.58 50.19 -49.04 50.65 ;
      RECT  -48.58 100.59 -49.04 101.05 ;
      RECT  -41.72 66.99 -42.18 67.45 ;
      RECT  -41.72 83.79 -42.18 84.25 ;
      RECT  -48.58 83.79 -49.04 84.25 ;
      RECT  -41.72 83.79 -42.18 84.25 ;
      RECT  -41.72 33.39 -42.18 33.85 ;
      RECT  -48.58 83.79 -49.04 84.25 ;
      RECT  -41.72 100.59 -42.18 101.05 ;
      RECT  -41.72 50.19 -42.18 50.65 ;
      RECT  -48.58 66.99 -49.04 67.45 ;
      RECT  -48.58 33.39 -49.04 33.85 ;
      RECT  -41.72 58.59 -42.18 59.05 ;
      RECT  -41.72 41.79 -42.18 42.25 ;
      RECT  -41.72 75.39 -42.18 75.85 ;
      RECT  -48.58 75.39 -49.04 75.85 ;
      RECT  -41.72 92.19 -42.18 92.65 ;
      RECT  -48.58 24.99 -49.04 25.45 ;
      RECT  -41.72 24.99 -42.18 25.45 ;
      RECT  -48.58 41.79 -49.04 42.25 ;
      RECT  -48.58 58.59 -49.04 59.05 ;
      RECT  -48.58 92.19 -49.04 92.65 ;
      RECT  -49.04 66.99 -48.58 67.45 ;
      RECT  -49.04 33.39 -48.58 33.85 ;
      RECT  -42.18 33.39 -41.72 33.85 ;
      RECT  -42.18 100.59 -41.72 101.05 ;
      RECT  -49.04 83.79 -48.58 84.25 ;
      RECT  -49.04 100.59 -48.58 101.05 ;
      RECT  -49.04 50.19 -48.58 50.65 ;
      RECT  -53.07 -6.02 -52.61 -5.56 ;
      RECT  -42.18 66.99 -41.72 67.45 ;
      RECT  -42.18 83.79 -41.72 84.25 ;
      RECT  -42.18 50.19 -41.72 50.65 ;
      RECT  -53.07 -6.04 -52.61 -5.58 ;
      RECT  -42.18 24.99 -41.72 25.45 ;
      RECT  -42.18 58.59 -41.72 59.05 ;
      RECT  -53.07 -1.8 -52.61 -1.34 ;
      RECT  -53.07 -10.26 -52.61 -9.8 ;
      RECT  -49.04 41.79 -48.58 42.25 ;
      RECT  -42.18 92.19 -41.72 92.65 ;
      RECT  -49.04 24.99 -48.58 25.45 ;
      RECT  -49.04 75.39 -48.58 75.85 ;
      RECT  -49.04 58.59 -48.58 59.05 ;
      RECT  -49.04 92.19 -48.58 92.65 ;
      RECT  -42.18 41.79 -41.72 42.25 ;
      RECT  -42.18 75.39 -41.72 75.85 ;
      RECT  -14.53 103.99 -1.4 104.29 ;
      RECT  -8.19 106.06 -7.73 106.52 ;
      RECT  -8.19 106.04 -7.73 106.5 ;
      RECT  -8.19 114.58 -7.73 115.04 ;
      RECT  -8.19 114.56 -7.73 115.02 ;
      RECT  -8.19 118.82 -7.73 119.28 ;
      RECT  -8.19 110.3 -7.73 110.76 ;
      RECT  -8.19 101.8 -7.73 102.26 ;
      RECT  -8.19 110.32 -7.73 110.78 ;
      RECT  11.73 -8.09 37.99 -7.79 ;
      RECT  18.07 -6.02 18.53 -5.56 ;
      RECT  31.19 -6.02 31.65 -5.56 ;
      RECT  18.07 -10.28 18.53 -9.82 ;
      RECT  31.19 -10.28 31.65 -9.82 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130A
END    LIBRARY
