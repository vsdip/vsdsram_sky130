magic
tech sky130A
timestamp 1616661915
<< nwell >>
rect 0 287 400 490
<< nmos >>
rect 78 210 93 252
rect 119 48 134 148
rect 241 48 256 90
rect 292 48 307 90
<< pmos >>
rect 78 333 93 388
rect 202 305 217 405
rect 292 305 307 360
<< ndiff >>
rect 38 240 78 252
rect 38 223 48 240
rect 65 223 78 240
rect 38 210 78 223
rect 93 240 138 252
rect 93 223 108 240
rect 125 223 138 240
rect 93 210 138 223
rect 79 78 119 148
rect 79 61 89 78
rect 106 61 119 78
rect 79 48 119 61
rect 134 121 179 148
rect 134 104 149 121
rect 166 104 179 121
rect 134 78 179 104
rect 134 61 149 78
rect 166 61 179 78
rect 134 48 179 61
rect 206 78 241 90
rect 206 61 214 78
rect 231 61 241 78
rect 206 48 241 61
rect 256 78 292 90
rect 256 61 266 78
rect 283 61 292 78
rect 256 48 292 61
rect 307 78 341 90
rect 307 61 316 78
rect 333 61 341 78
rect 307 48 341 61
<< pdiff >>
rect 165 394 202 405
rect 38 369 78 388
rect 38 352 48 369
rect 65 352 78 369
rect 38 333 78 352
rect 93 369 138 388
rect 93 352 108 369
rect 125 352 138 369
rect 93 333 138 352
rect 165 377 175 394
rect 192 377 202 394
rect 165 341 202 377
rect 165 324 175 341
rect 192 324 202 341
rect 165 305 202 324
rect 217 394 256 405
rect 217 377 226 394
rect 243 377 256 394
rect 217 360 256 377
rect 217 341 292 360
rect 217 324 226 341
rect 243 324 266 341
rect 283 324 292 341
rect 217 305 292 324
rect 307 341 341 360
rect 307 324 316 341
rect 333 324 341 341
rect 307 305 341 324
<< ndiffc >>
rect 48 223 65 240
rect 108 223 125 240
rect 89 61 106 78
rect 149 104 166 121
rect 149 61 166 78
rect 214 61 231 78
rect 266 61 283 78
rect 316 61 333 78
<< pdiffc >>
rect 48 352 65 369
rect 108 352 125 369
rect 175 377 192 394
rect 175 324 192 341
rect 226 377 243 394
rect 226 324 243 341
rect 266 324 283 341
rect 316 324 333 341
<< psubdiff >>
rect 79 8 120 20
rect 79 -9 91 8
rect 108 -9 120 8
rect 79 -21 120 -9
rect 248 8 289 20
rect 248 -9 260 8
rect 277 -9 289 8
rect 248 -21 289 -9
<< nsubdiff >>
rect 57 454 110 472
rect 57 437 75 454
rect 92 437 110 454
rect 57 419 110 437
<< psubdiffcont >>
rect 91 -9 108 8
rect 260 -9 277 8
<< nsubdiffcont >>
rect 75 437 92 454
<< poly >>
rect 202 405 217 422
rect 78 388 93 405
rect 78 299 93 333
rect 292 360 307 377
rect 78 291 117 299
rect 78 274 92 291
rect 109 274 117 291
rect 202 297 217 305
rect 292 297 307 305
rect 202 279 307 297
rect 78 266 117 274
rect 78 252 93 266
rect 150 221 183 229
rect 280 222 295 279
rect 78 195 93 210
rect 150 204 158 221
rect 175 220 183 221
rect 175 204 241 220
rect 150 196 183 204
rect 24 178 57 186
rect 24 161 32 178
rect 49 173 57 178
rect 49 161 134 173
rect 24 158 134 161
rect 24 153 57 158
rect 119 148 134 158
rect 226 113 241 204
rect 273 214 306 222
rect 273 197 281 214
rect 298 197 306 214
rect 273 189 306 197
rect 274 159 307 167
rect 274 142 282 159
rect 299 142 307 159
rect 274 134 307 142
rect 226 98 256 113
rect 241 90 256 98
rect 292 90 307 134
rect 119 33 134 48
rect 241 33 256 48
rect 292 33 307 48
<< polycont >>
rect 92 274 109 291
rect 158 204 175 221
rect 32 161 49 178
rect 281 197 298 214
rect 282 142 299 159
<< locali >>
rect 67 454 100 462
rect 0 437 75 454
rect 92 437 330 454
rect 347 437 400 454
rect 67 429 117 437
rect 100 377 117 429
rect 218 402 237 437
rect 167 394 200 402
rect 167 377 175 394
rect 192 377 200 394
rect 40 369 73 377
rect 40 352 48 369
rect 65 352 73 369
rect 40 344 73 352
rect 100 369 133 377
rect 100 352 108 369
rect 125 352 133 369
rect 100 344 133 352
rect 48 315 65 344
rect 167 341 200 377
rect 167 324 175 341
rect 192 324 200 341
rect 167 316 200 324
rect 218 394 251 402
rect 218 377 226 394
rect 243 377 251 394
rect 218 349 251 377
rect 218 341 291 349
rect 218 324 226 341
rect 243 324 266 341
rect 283 324 291 341
rect 218 316 291 324
rect 308 341 341 349
rect 308 324 316 341
rect 333 324 341 341
rect 308 316 341 324
rect 59 298 65 315
rect 48 248 65 298
rect 84 291 117 299
rect 173 291 190 316
rect 84 274 92 291
rect 109 275 190 291
rect 109 274 239 275
rect 84 266 117 274
rect 173 258 239 274
rect 40 240 73 248
rect 40 223 48 240
rect 65 223 73 240
rect 40 215 73 223
rect 100 240 133 248
rect 100 223 108 240
rect 125 223 133 240
rect 100 215 133 223
rect 150 221 183 229
rect 114 191 131 215
rect 150 204 158 221
rect 175 204 183 221
rect 150 196 183 204
rect 24 178 57 186
rect 24 161 32 178
rect 49 161 57 178
rect 24 153 57 161
rect 81 174 131 191
rect 81 89 98 174
rect 141 121 174 129
rect 141 104 149 121
rect 166 104 174 121
rect 81 78 114 89
rect 81 61 89 78
rect 106 61 114 78
rect 81 53 114 61
rect 141 78 174 104
rect 222 86 239 258
rect 273 220 306 222
rect 324 220 341 316
rect 273 214 341 220
rect 273 197 281 214
rect 298 203 341 214
rect 298 197 306 203
rect 273 189 306 197
rect 274 159 307 167
rect 274 142 282 159
rect 299 142 307 159
rect 274 134 307 142
rect 141 61 149 78
rect 166 61 174 78
rect 141 53 174 61
rect 198 78 239 86
rect 198 61 214 78
rect 231 61 239 78
rect 198 53 239 61
rect 258 78 291 86
rect 324 83 341 203
rect 258 61 266 78
rect 283 61 291 78
rect 258 53 291 61
rect 308 78 341 83
rect 308 61 316 78
rect 333 61 341 78
rect 308 53 341 61
rect 91 16 108 53
rect 83 8 116 16
rect 252 8 285 16
rect 0 -9 91 8
rect 108 -9 153 8
rect 170 -9 260 8
rect 277 -9 345 8
rect 362 -9 400 8
rect 83 -17 116 -9
rect 252 -17 285 -9
<< viali >>
rect 75 437 92 454
rect 330 437 347 454
rect 42 298 59 315
rect 158 204 175 221
rect 32 161 49 178
rect 282 142 299 159
rect 149 61 166 78
rect 266 61 283 78
rect 91 -9 108 8
rect 153 -9 170 8
rect 260 -9 277 8
rect 345 -9 362 8
<< metal1 >>
rect 0 454 324 460
rect 0 437 75 454
rect 92 437 324 454
rect 0 431 324 437
rect 353 431 400 460
rect 36 315 65 321
rect 36 312 42 315
rect 0 298 42 312
rect 59 312 65 315
rect 59 298 400 312
rect 36 292 65 298
rect 150 225 183 229
rect 150 199 153 225
rect 179 199 183 225
rect 150 196 183 199
rect 26 179 55 184
rect 26 178 57 179
rect 26 161 32 178
rect 49 161 57 178
rect 26 155 57 161
rect 43 113 57 155
rect 274 163 307 167
rect 274 137 277 163
rect 303 137 307 163
rect 274 134 307 137
rect 0 99 400 113
rect 143 78 172 84
rect 143 61 149 78
rect 166 75 172 78
rect 260 78 289 84
rect 260 75 266 78
rect 166 61 266 75
rect 283 61 289 78
rect 143 55 172 61
rect 260 55 289 61
rect 0 8 338 14
rect 0 -9 91 8
rect 108 -9 153 8
rect 170 -9 260 8
rect 277 -9 338 8
rect 0 -15 338 -9
rect 367 -15 400 14
<< via1 >>
rect 324 454 353 460
rect 324 437 330 454
rect 330 437 347 454
rect 347 437 353 454
rect 324 431 353 437
rect 153 221 179 225
rect 153 204 158 221
rect 158 204 175 221
rect 175 204 179 221
rect 153 199 179 204
rect 277 159 303 163
rect 277 142 282 159
rect 282 142 299 159
rect 299 142 303 159
rect 277 137 303 142
rect 338 8 367 14
rect 338 -9 345 8
rect 345 -9 362 8
rect 362 -9 367 8
rect 338 -15 367 -9
<< metal2 >>
rect 150 229 164 490
rect 150 225 183 229
rect 150 199 153 225
rect 179 199 183 225
rect 150 196 183 199
rect 150 -21 164 196
rect 261 167 275 490
rect 316 463 361 468
rect 316 428 321 463
rect 356 428 361 463
rect 316 423 361 428
rect 261 163 307 167
rect 261 137 277 163
rect 303 137 307 163
rect 261 134 307 137
rect 261 -21 275 134
rect 330 17 375 22
rect 330 -18 335 17
rect 370 -18 375 17
rect 330 -23 375 -18
<< via2 >>
rect 321 460 356 463
rect 321 431 324 460
rect 324 431 353 460
rect 353 431 356 460
rect 321 428 356 431
rect 335 14 370 17
rect 335 -15 338 14
rect 338 -15 367 14
rect 367 -15 370 14
rect 335 -18 370 -15
<< metal3 >>
rect 310 463 363 470
rect 310 428 321 463
rect 356 428 363 463
rect 310 420 363 428
rect 325 17 377 25
rect 325 -18 335 17
rect 370 -18 377 17
rect 325 -25 377 -18
<< labels >>
flabel metal1 s 44 301 58 314 0 FreeSans 200 180 0 0 dout
port 17 nsew
flabel metal1 s 170 -5 183 5 0 FreeSans 200 180 0 0 gnd
port 20 nsew
flabel metal2 s 285 144 297 157 0 FreeSans 200 180 0 0 br
port 16 nsew
flabel metal1 s 34 160 48 173 0 FreeSans 200 180 0 0 en
port 18 nsew
flabel metal1 s 217 440 230 450 0 FreeSans 200 180 0 0 vdd
port 19 nsew
flabel metal2 s 161 207 173 219 0 FreeSans 200 180 0 0 bl
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 400 445
<< end >>
